module r_ram_for_sign
(
	input wire clk,
	input wire reset,
    input r_ram_for_sign_start,
	input [7:0] data, 


	output[14:0] address,
    output [19584-1:0] sigma_out,
	output reg  r_ram_for_sign_end
);


// M 6399
reg [7:0]M_list[6399:0];
wire [51199:0]M={M_list[0],M_list[1],M_list[2],M_list[3],M_list[4],M_list[5],M_list[6],M_list[7],M_list[8],M_list[9],M_list[10],M_list[11],M_list[12],M_list[13],M_list[14],M_list[15],M_list[16],M_list[17],M_list[18],M_list[19],M_list[20],M_list[21],M_list[22],M_list[23],M_list[24],M_list[25],M_list[26],M_list[27],M_list[28],M_list[29],M_list[30],M_list[31],M_list[32],M_list[33],M_list[34],M_list[35],M_list[36],M_list[37],M_list[38],M_list[39],M_list[40],M_list[41],M_list[42],M_list[43],M_list[44],M_list[45],M_list[46],M_list[47],M_list[48],M_list[49],M_list[50],M_list[51],M_list[52],M_list[53],M_list[54],M_list[55],M_list[56],M_list[57],M_list[58],M_list[59],M_list[60],M_list[61],M_list[62],M_list[63],M_list[64],M_list[65],M_list[66],M_list[67],M_list[68],M_list[69],M_list[70],M_list[71],M_list[72],M_list[73],M_list[74],M_list[75],M_list[76],M_list[77],M_list[78],M_list[79],M_list[80],M_list[81],M_list[82],M_list[83],M_list[84],M_list[85],M_list[86],M_list[87],M_list[88],M_list[89],M_list[90],M_list[91],M_list[92],M_list[93],M_list[94],M_list[95],M_list[96],M_list[97],M_list[98],M_list[99],M_list[100],M_list[101],M_list[102],M_list[103],M_list[104],M_list[105],M_list[106],M_list[107],M_list[108],M_list[109],M_list[110],M_list[111],M_list[112],M_list[113],M_list[114],M_list[115],M_list[116],M_list[117],M_list[118],M_list[119],M_list[120],M_list[121],M_list[122],M_list[123],M_list[124],M_list[125],M_list[126],M_list[127],M_list[128],M_list[129],M_list[130],M_list[131],M_list[132],M_list[133],M_list[134],M_list[135],M_list[136],M_list[137],M_list[138],M_list[139],M_list[140],M_list[141],M_list[142],M_list[143],M_list[144],M_list[145],M_list[146],M_list[147],M_list[148],M_list[149],M_list[150],M_list[151],M_list[152],M_list[153],M_list[154],M_list[155],M_list[156],M_list[157],M_list[158],M_list[159],M_list[160],M_list[161],M_list[162],M_list[163],M_list[164],M_list[165],M_list[166],M_list[167],M_list[168],M_list[169],M_list[170],M_list[171],M_list[172],M_list[173],M_list[174],M_list[175],M_list[176],M_list[177],M_list[178],M_list[179],M_list[180],M_list[181],M_list[182],M_list[183],M_list[184],M_list[185],M_list[186],M_list[187],M_list[188],M_list[189],M_list[190],M_list[191],M_list[192],M_list[193],M_list[194],M_list[195],M_list[196],M_list[197],M_list[198],M_list[199],M_list[200],M_list[201],M_list[202],M_list[203],M_list[204],M_list[205],M_list[206],M_list[207],M_list[208],M_list[209],M_list[210],M_list[211],M_list[212],M_list[213],M_list[214],M_list[215],M_list[216],M_list[217],M_list[218],M_list[219],M_list[220],M_list[221],M_list[222],M_list[223],M_list[224],M_list[225],M_list[226],M_list[227],M_list[228],M_list[229],M_list[230],M_list[231],M_list[232],M_list[233],M_list[234],M_list[235],M_list[236],M_list[237],M_list[238],M_list[239],M_list[240],M_list[241],M_list[242],M_list[243],M_list[244],M_list[245],M_list[246],M_list[247],M_list[248],M_list[249],M_list[250],M_list[251],M_list[252],M_list[253],M_list[254],M_list[255],M_list[256],M_list[257],M_list[258],M_list[259],M_list[260],M_list[261],M_list[262],M_list[263],M_list[264],M_list[265],M_list[266],M_list[267],M_list[268],M_list[269],M_list[270],M_list[271],M_list[272],M_list[273],M_list[274],M_list[275],M_list[276],M_list[277],M_list[278],M_list[279],M_list[280],M_list[281],M_list[282],M_list[283],M_list[284],M_list[285],M_list[286],M_list[287],M_list[288],M_list[289],M_list[290],M_list[291],M_list[292],M_list[293],M_list[294],M_list[295],M_list[296],M_list[297],M_list[298],M_list[299],M_list[300],M_list[301],M_list[302],M_list[303],M_list[304],M_list[305],M_list[306],M_list[307],M_list[308],M_list[309],M_list[310],M_list[311],M_list[312],M_list[313],M_list[314],M_list[315],M_list[316],M_list[317],M_list[318],M_list[319],M_list[320],M_list[321],M_list[322],M_list[323],M_list[324],M_list[325],M_list[326],M_list[327],M_list[328],M_list[329],M_list[330],M_list[331],M_list[332],M_list[333],M_list[334],M_list[335],M_list[336],M_list[337],M_list[338],M_list[339],M_list[340],M_list[341],M_list[342],M_list[343],M_list[344],M_list[345],M_list[346],M_list[347],M_list[348],M_list[349],M_list[350],M_list[351],M_list[352],M_list[353],M_list[354],M_list[355],M_list[356],M_list[357],M_list[358],M_list[359],M_list[360],M_list[361],M_list[362],M_list[363],M_list[364],M_list[365],M_list[366],M_list[367],M_list[368],M_list[369],M_list[370],M_list[371],M_list[372],M_list[373],M_list[374],M_list[375],M_list[376],M_list[377],M_list[378],M_list[379],M_list[380],M_list[381],M_list[382],M_list[383],M_list[384],M_list[385],M_list[386],M_list[387],M_list[388],M_list[389],M_list[390],M_list[391],M_list[392],M_list[393],M_list[394],M_list[395],M_list[396],M_list[397],M_list[398],M_list[399],M_list[400],M_list[401],M_list[402],M_list[403],M_list[404],M_list[405],M_list[406],M_list[407],M_list[408],M_list[409],M_list[410],M_list[411],M_list[412],M_list[413],M_list[414],M_list[415],M_list[416],M_list[417],M_list[418],M_list[419],M_list[420],M_list[421],M_list[422],M_list[423],M_list[424],M_list[425],M_list[426],M_list[427],M_list[428],M_list[429],M_list[430],M_list[431],M_list[432],M_list[433],M_list[434],M_list[435],M_list[436],M_list[437],M_list[438],M_list[439],M_list[440],M_list[441],M_list[442],M_list[443],M_list[444],M_list[445],M_list[446],M_list[447],M_list[448],M_list[449],M_list[450],M_list[451],M_list[452],M_list[453],M_list[454],M_list[455],M_list[456],M_list[457],M_list[458],M_list[459],M_list[460],M_list[461],M_list[462],M_list[463],M_list[464],M_list[465],M_list[466],M_list[467],M_list[468],M_list[469],M_list[470],M_list[471],M_list[472],M_list[473],M_list[474],M_list[475],M_list[476],M_list[477],M_list[478],M_list[479],M_list[480],M_list[481],M_list[482],M_list[483],M_list[484],M_list[485],M_list[486],M_list[487],M_list[488],M_list[489],M_list[490],M_list[491],M_list[492],M_list[493],M_list[494],M_list[495],M_list[496],M_list[497],M_list[498],M_list[499],M_list[500],M_list[501],M_list[502],M_list[503],M_list[504],M_list[505],M_list[506],M_list[507],M_list[508],M_list[509],M_list[510],M_list[511],M_list[512],M_list[513],M_list[514],M_list[515],M_list[516],M_list[517],M_list[518],M_list[519],M_list[520],M_list[521],M_list[522],M_list[523],M_list[524],M_list[525],M_list[526],M_list[527],M_list[528],M_list[529],M_list[530],M_list[531],M_list[532],M_list[533],M_list[534],M_list[535],M_list[536],M_list[537],M_list[538],M_list[539],M_list[540],M_list[541],M_list[542],M_list[543],M_list[544],M_list[545],M_list[546],M_list[547],M_list[548],M_list[549],M_list[550],M_list[551],M_list[552],M_list[553],M_list[554],M_list[555],M_list[556],M_list[557],M_list[558],M_list[559],M_list[560],M_list[561],M_list[562],M_list[563],M_list[564],M_list[565],M_list[566],M_list[567],M_list[568],M_list[569],M_list[570],M_list[571],M_list[572],M_list[573],M_list[574],M_list[575],M_list[576],M_list[577],M_list[578],M_list[579],M_list[580],M_list[581],M_list[582],M_list[583],M_list[584],M_list[585],M_list[586],M_list[587],M_list[588],M_list[589],M_list[590],M_list[591],M_list[592],M_list[593],M_list[594],M_list[595],M_list[596],M_list[597],M_list[598],M_list[599],M_list[600],M_list[601],M_list[602],M_list[603],M_list[604],M_list[605],M_list[606],M_list[607],M_list[608],M_list[609],M_list[610],M_list[611],M_list[612],M_list[613],M_list[614],M_list[615],M_list[616],M_list[617],M_list[618],M_list[619],M_list[620],M_list[621],M_list[622],M_list[623],M_list[624],M_list[625],M_list[626],M_list[627],M_list[628],M_list[629],M_list[630],M_list[631],M_list[632],M_list[633],M_list[634],M_list[635],M_list[636],M_list[637],M_list[638],M_list[639],M_list[640],M_list[641],M_list[642],M_list[643],M_list[644],M_list[645],M_list[646],M_list[647],M_list[648],M_list[649],M_list[650],M_list[651],M_list[652],M_list[653],M_list[654],M_list[655],M_list[656],M_list[657],M_list[658],M_list[659],M_list[660],M_list[661],M_list[662],M_list[663],M_list[664],M_list[665],M_list[666],M_list[667],M_list[668],M_list[669],M_list[670],M_list[671],M_list[672],M_list[673],M_list[674],M_list[675],M_list[676],M_list[677],M_list[678],M_list[679],M_list[680],M_list[681],M_list[682],M_list[683],M_list[684],M_list[685],M_list[686],M_list[687],M_list[688],M_list[689],M_list[690],M_list[691],M_list[692],M_list[693],M_list[694],M_list[695],M_list[696],M_list[697],M_list[698],M_list[699],M_list[700],M_list[701],M_list[702],M_list[703],M_list[704],M_list[705],M_list[706],M_list[707],M_list[708],M_list[709],M_list[710],M_list[711],M_list[712],M_list[713],M_list[714],M_list[715],M_list[716],M_list[717],M_list[718],M_list[719],M_list[720],M_list[721],M_list[722],M_list[723],M_list[724],M_list[725],M_list[726],M_list[727],M_list[728],M_list[729],M_list[730],M_list[731],M_list[732],M_list[733],M_list[734],M_list[735],M_list[736],M_list[737],M_list[738],M_list[739],M_list[740],M_list[741],M_list[742],M_list[743],M_list[744],M_list[745],M_list[746],M_list[747],M_list[748],M_list[749],M_list[750],M_list[751],M_list[752],M_list[753],M_list[754],M_list[755],M_list[756],M_list[757],M_list[758],M_list[759],M_list[760],M_list[761],M_list[762],M_list[763],M_list[764],M_list[765],M_list[766],M_list[767],M_list[768],M_list[769],M_list[770],M_list[771],M_list[772],M_list[773],M_list[774],M_list[775],M_list[776],M_list[777],M_list[778],M_list[779],M_list[780],M_list[781],M_list[782],M_list[783],M_list[784],M_list[785],M_list[786],M_list[787],M_list[788],M_list[789],M_list[790],M_list[791],M_list[792],M_list[793],M_list[794],M_list[795],M_list[796],M_list[797],M_list[798],M_list[799],M_list[800],M_list[801],M_list[802],M_list[803],M_list[804],M_list[805],M_list[806],M_list[807],M_list[808],M_list[809],M_list[810],M_list[811],M_list[812],M_list[813],M_list[814],M_list[815],M_list[816],M_list[817],M_list[818],M_list[819],M_list[820],M_list[821],M_list[822],M_list[823],M_list[824],M_list[825],M_list[826],M_list[827],M_list[828],M_list[829],M_list[830],M_list[831],M_list[832],M_list[833],M_list[834],M_list[835],M_list[836],M_list[837],M_list[838],M_list[839],M_list[840],M_list[841],M_list[842],M_list[843],M_list[844],M_list[845],M_list[846],M_list[847],M_list[848],M_list[849],M_list[850],M_list[851],M_list[852],M_list[853],M_list[854],M_list[855],M_list[856],M_list[857],M_list[858],M_list[859],M_list[860],M_list[861],M_list[862],M_list[863],M_list[864],M_list[865],M_list[866],M_list[867],M_list[868],M_list[869],M_list[870],M_list[871],M_list[872],M_list[873],M_list[874],M_list[875],M_list[876],M_list[877],M_list[878],M_list[879],M_list[880],M_list[881],M_list[882],M_list[883],M_list[884],M_list[885],M_list[886],M_list[887],M_list[888],M_list[889],M_list[890],M_list[891],M_list[892],M_list[893],M_list[894],M_list[895],M_list[896],M_list[897],M_list[898],M_list[899],M_list[900],M_list[901],M_list[902],M_list[903],M_list[904],M_list[905],M_list[906],M_list[907],M_list[908],M_list[909],M_list[910],M_list[911],M_list[912],M_list[913],M_list[914],M_list[915],M_list[916],M_list[917],M_list[918],M_list[919],M_list[920],M_list[921],M_list[922],M_list[923],M_list[924],M_list[925],M_list[926],M_list[927],M_list[928],M_list[929],M_list[930],M_list[931],M_list[932],M_list[933],M_list[934],M_list[935],M_list[936],M_list[937],M_list[938],M_list[939],M_list[940],M_list[941],M_list[942],M_list[943],M_list[944],M_list[945],M_list[946],M_list[947],M_list[948],M_list[949],M_list[950],M_list[951],M_list[952],M_list[953],M_list[954],M_list[955],M_list[956],M_list[957],M_list[958],M_list[959],M_list[960],M_list[961],M_list[962],M_list[963],M_list[964],M_list[965],M_list[966],M_list[967],M_list[968],M_list[969],M_list[970],M_list[971],M_list[972],M_list[973],M_list[974],M_list[975],M_list[976],M_list[977],M_list[978],M_list[979],M_list[980],M_list[981],M_list[982],M_list[983],M_list[984],M_list[985],M_list[986],M_list[987],M_list[988],M_list[989],M_list[990],M_list[991],M_list[992],M_list[993],M_list[994],M_list[995],M_list[996],M_list[997],M_list[998],M_list[999],M_list[1000],M_list[1001],M_list[1002],M_list[1003],M_list[1004],M_list[1005],M_list[1006],M_list[1007],M_list[1008],M_list[1009],M_list[1010],M_list[1011],M_list[1012],M_list[1013],M_list[1014],M_list[1015],M_list[1016],M_list[1017],M_list[1018],M_list[1019],M_list[1020],M_list[1021],M_list[1022],M_list[1023],M_list[1024],M_list[1025],M_list[1026],M_list[1027],M_list[1028],M_list[1029],M_list[1030],M_list[1031],M_list[1032],M_list[1033],M_list[1034],M_list[1035],M_list[1036],M_list[1037],M_list[1038],M_list[1039],M_list[1040],M_list[1041],M_list[1042],M_list[1043],M_list[1044],M_list[1045],M_list[1046],M_list[1047],M_list[1048],M_list[1049],M_list[1050],M_list[1051],M_list[1052],M_list[1053],M_list[1054],M_list[1055],M_list[1056],M_list[1057],M_list[1058],M_list[1059],M_list[1060],M_list[1061],M_list[1062],M_list[1063],M_list[1064],M_list[1065],M_list[1066],M_list[1067],M_list[1068],M_list[1069],M_list[1070],M_list[1071],M_list[1072],M_list[1073],M_list[1074],M_list[1075],M_list[1076],M_list[1077],M_list[1078],M_list[1079],M_list[1080],M_list[1081],M_list[1082],M_list[1083],M_list[1084],M_list[1085],M_list[1086],M_list[1087],M_list[1088],M_list[1089],M_list[1090],M_list[1091],M_list[1092],M_list[1093],M_list[1094],M_list[1095],M_list[1096],M_list[1097],M_list[1098],M_list[1099],M_list[1100],M_list[1101],M_list[1102],M_list[1103],M_list[1104],M_list[1105],M_list[1106],M_list[1107],M_list[1108],M_list[1109],M_list[1110],M_list[1111],M_list[1112],M_list[1113],M_list[1114],M_list[1115],M_list[1116],M_list[1117],M_list[1118],M_list[1119],M_list[1120],M_list[1121],M_list[1122],M_list[1123],M_list[1124],M_list[1125],M_list[1126],M_list[1127],M_list[1128],M_list[1129],M_list[1130],M_list[1131],M_list[1132],M_list[1133],M_list[1134],M_list[1135],M_list[1136],M_list[1137],M_list[1138],M_list[1139],M_list[1140],M_list[1141],M_list[1142],M_list[1143],M_list[1144],M_list[1145],M_list[1146],M_list[1147],M_list[1148],M_list[1149],M_list[1150],M_list[1151],M_list[1152],M_list[1153],M_list[1154],M_list[1155],M_list[1156],M_list[1157],M_list[1158],M_list[1159],M_list[1160],M_list[1161],M_list[1162],M_list[1163],M_list[1164],M_list[1165],M_list[1166],M_list[1167],M_list[1168],M_list[1169],M_list[1170],M_list[1171],M_list[1172],M_list[1173],M_list[1174],M_list[1175],M_list[1176],M_list[1177],M_list[1178],M_list[1179],M_list[1180],M_list[1181],M_list[1182],M_list[1183],M_list[1184],M_list[1185],M_list[1186],M_list[1187],M_list[1188],M_list[1189],M_list[1190],M_list[1191],M_list[1192],M_list[1193],M_list[1194],M_list[1195],M_list[1196],M_list[1197],M_list[1198],M_list[1199],M_list[1200],M_list[1201],M_list[1202],M_list[1203],M_list[1204],M_list[1205],M_list[1206],M_list[1207],M_list[1208],M_list[1209],M_list[1210],M_list[1211],M_list[1212],M_list[1213],M_list[1214],M_list[1215],M_list[1216],M_list[1217],M_list[1218],M_list[1219],M_list[1220],M_list[1221],M_list[1222],M_list[1223],M_list[1224],M_list[1225],M_list[1226],M_list[1227],M_list[1228],M_list[1229],M_list[1230],M_list[1231],M_list[1232],M_list[1233],M_list[1234],M_list[1235],M_list[1236],M_list[1237],M_list[1238],M_list[1239],M_list[1240],M_list[1241],M_list[1242],M_list[1243],M_list[1244],M_list[1245],M_list[1246],M_list[1247],M_list[1248],M_list[1249],M_list[1250],M_list[1251],M_list[1252],M_list[1253],M_list[1254],M_list[1255],M_list[1256],M_list[1257],M_list[1258],M_list[1259],M_list[1260],M_list[1261],M_list[1262],M_list[1263],M_list[1264],M_list[1265],M_list[1266],M_list[1267],M_list[1268],M_list[1269],M_list[1270],M_list[1271],M_list[1272],M_list[1273],M_list[1274],M_list[1275],M_list[1276],M_list[1277],M_list[1278],M_list[1279],M_list[1280],M_list[1281],M_list[1282],M_list[1283],M_list[1284],M_list[1285],M_list[1286],M_list[1287],M_list[1288],M_list[1289],M_list[1290],M_list[1291],M_list[1292],M_list[1293],M_list[1294],M_list[1295],M_list[1296],M_list[1297],M_list[1298],M_list[1299],M_list[1300],M_list[1301],M_list[1302],M_list[1303],M_list[1304],M_list[1305],M_list[1306],M_list[1307],M_list[1308],M_list[1309],M_list[1310],M_list[1311],M_list[1312],M_list[1313],M_list[1314],M_list[1315],M_list[1316],M_list[1317],M_list[1318],M_list[1319],M_list[1320],M_list[1321],M_list[1322],M_list[1323],M_list[1324],M_list[1325],M_list[1326],M_list[1327],M_list[1328],M_list[1329],M_list[1330],M_list[1331],M_list[1332],M_list[1333],M_list[1334],M_list[1335],M_list[1336],M_list[1337],M_list[1338],M_list[1339],M_list[1340],M_list[1341],M_list[1342],M_list[1343],M_list[1344],M_list[1345],M_list[1346],M_list[1347],M_list[1348],M_list[1349],M_list[1350],M_list[1351],M_list[1352],M_list[1353],M_list[1354],M_list[1355],M_list[1356],M_list[1357],M_list[1358],M_list[1359],M_list[1360],M_list[1361],M_list[1362],M_list[1363],M_list[1364],M_list[1365],M_list[1366],M_list[1367],M_list[1368],M_list[1369],M_list[1370],M_list[1371],M_list[1372],M_list[1373],M_list[1374],M_list[1375],M_list[1376],M_list[1377],M_list[1378],M_list[1379],M_list[1380],M_list[1381],M_list[1382],M_list[1383],M_list[1384],M_list[1385],M_list[1386],M_list[1387],M_list[1388],M_list[1389],M_list[1390],M_list[1391],M_list[1392],M_list[1393],M_list[1394],M_list[1395],M_list[1396],M_list[1397],M_list[1398],M_list[1399],M_list[1400],M_list[1401],M_list[1402],M_list[1403],M_list[1404],M_list[1405],M_list[1406],M_list[1407],M_list[1408],M_list[1409],M_list[1410],M_list[1411],M_list[1412],M_list[1413],M_list[1414],M_list[1415],M_list[1416],M_list[1417],M_list[1418],M_list[1419],M_list[1420],M_list[1421],M_list[1422],M_list[1423],M_list[1424],M_list[1425],M_list[1426],M_list[1427],M_list[1428],M_list[1429],M_list[1430],M_list[1431],M_list[1432],M_list[1433],M_list[1434],M_list[1435],M_list[1436],M_list[1437],M_list[1438],M_list[1439],M_list[1440],M_list[1441],M_list[1442],M_list[1443],M_list[1444],M_list[1445],M_list[1446],M_list[1447],M_list[1448],M_list[1449],M_list[1450],M_list[1451],M_list[1452],M_list[1453],M_list[1454],M_list[1455],M_list[1456],M_list[1457],M_list[1458],M_list[1459],M_list[1460],M_list[1461],M_list[1462],M_list[1463],M_list[1464],M_list[1465],M_list[1466],M_list[1467],M_list[1468],M_list[1469],M_list[1470],M_list[1471],M_list[1472],M_list[1473],M_list[1474],M_list[1475],M_list[1476],M_list[1477],M_list[1478],M_list[1479],M_list[1480],M_list[1481],M_list[1482],M_list[1483],M_list[1484],M_list[1485],M_list[1486],M_list[1487],M_list[1488],M_list[1489],M_list[1490],M_list[1491],M_list[1492],M_list[1493],M_list[1494],M_list[1495],M_list[1496],M_list[1497],M_list[1498],M_list[1499],M_list[1500],M_list[1501],M_list[1502],M_list[1503],M_list[1504],M_list[1505],M_list[1506],M_list[1507],M_list[1508],M_list[1509],M_list[1510],M_list[1511],M_list[1512],M_list[1513],M_list[1514],M_list[1515],M_list[1516],M_list[1517],M_list[1518],M_list[1519],M_list[1520],M_list[1521],M_list[1522],M_list[1523],M_list[1524],M_list[1525],M_list[1526],M_list[1527],M_list[1528],M_list[1529],M_list[1530],M_list[1531],M_list[1532],M_list[1533],M_list[1534],M_list[1535],M_list[1536],M_list[1537],M_list[1538],M_list[1539],M_list[1540],M_list[1541],M_list[1542],M_list[1543],M_list[1544],M_list[1545],M_list[1546],M_list[1547],M_list[1548],M_list[1549],M_list[1550],M_list[1551],M_list[1552],M_list[1553],M_list[1554],M_list[1555],M_list[1556],M_list[1557],M_list[1558],M_list[1559],M_list[1560],M_list[1561],M_list[1562],M_list[1563],M_list[1564],M_list[1565],M_list[1566],M_list[1567],M_list[1568],M_list[1569],M_list[1570],M_list[1571],M_list[1572],M_list[1573],M_list[1574],M_list[1575],M_list[1576],M_list[1577],M_list[1578],M_list[1579],M_list[1580],M_list[1581],M_list[1582],M_list[1583],M_list[1584],M_list[1585],M_list[1586],M_list[1587],M_list[1588],M_list[1589],M_list[1590],M_list[1591],M_list[1592],M_list[1593],M_list[1594],M_list[1595],M_list[1596],M_list[1597],M_list[1598],M_list[1599],M_list[1600],M_list[1601],M_list[1602],M_list[1603],M_list[1604],M_list[1605],M_list[1606],M_list[1607],M_list[1608],M_list[1609],M_list[1610],M_list[1611],M_list[1612],M_list[1613],M_list[1614],M_list[1615],M_list[1616],M_list[1617],M_list[1618],M_list[1619],M_list[1620],M_list[1621],M_list[1622],M_list[1623],M_list[1624],M_list[1625],M_list[1626],M_list[1627],M_list[1628],M_list[1629],M_list[1630],M_list[1631],M_list[1632],M_list[1633],M_list[1634],M_list[1635],M_list[1636],M_list[1637],M_list[1638],M_list[1639],M_list[1640],M_list[1641],M_list[1642],M_list[1643],M_list[1644],M_list[1645],M_list[1646],M_list[1647],M_list[1648],M_list[1649],M_list[1650],M_list[1651],M_list[1652],M_list[1653],M_list[1654],M_list[1655],M_list[1656],M_list[1657],M_list[1658],M_list[1659],M_list[1660],M_list[1661],M_list[1662],M_list[1663],M_list[1664],M_list[1665],M_list[1666],M_list[1667],M_list[1668],M_list[1669],M_list[1670],M_list[1671],M_list[1672],M_list[1673],M_list[1674],M_list[1675],M_list[1676],M_list[1677],M_list[1678],M_list[1679],M_list[1680],M_list[1681],M_list[1682],M_list[1683],M_list[1684],M_list[1685],M_list[1686],M_list[1687],M_list[1688],M_list[1689],M_list[1690],M_list[1691],M_list[1692],M_list[1693],M_list[1694],M_list[1695],M_list[1696],M_list[1697],M_list[1698],M_list[1699],M_list[1700],M_list[1701],M_list[1702],M_list[1703],M_list[1704],M_list[1705],M_list[1706],M_list[1707],M_list[1708],M_list[1709],M_list[1710],M_list[1711],M_list[1712],M_list[1713],M_list[1714],M_list[1715],M_list[1716],M_list[1717],M_list[1718],M_list[1719],M_list[1720],M_list[1721],M_list[1722],M_list[1723],M_list[1724],M_list[1725],M_list[1726],M_list[1727],M_list[1728],M_list[1729],M_list[1730],M_list[1731],M_list[1732],M_list[1733],M_list[1734],M_list[1735],M_list[1736],M_list[1737],M_list[1738],M_list[1739],M_list[1740],M_list[1741],M_list[1742],M_list[1743],M_list[1744],M_list[1745],M_list[1746],M_list[1747],M_list[1748],M_list[1749],M_list[1750],M_list[1751],M_list[1752],M_list[1753],M_list[1754],M_list[1755],M_list[1756],M_list[1757],M_list[1758],M_list[1759],M_list[1760],M_list[1761],M_list[1762],M_list[1763],M_list[1764],M_list[1765],M_list[1766],M_list[1767],M_list[1768],M_list[1769],M_list[1770],M_list[1771],M_list[1772],M_list[1773],M_list[1774],M_list[1775],M_list[1776],M_list[1777],M_list[1778],M_list[1779],M_list[1780],M_list[1781],M_list[1782],M_list[1783],M_list[1784],M_list[1785],M_list[1786],M_list[1787],M_list[1788],M_list[1789],M_list[1790],M_list[1791],M_list[1792],M_list[1793],M_list[1794],M_list[1795],M_list[1796],M_list[1797],M_list[1798],M_list[1799],M_list[1800],M_list[1801],M_list[1802],M_list[1803],M_list[1804],M_list[1805],M_list[1806],M_list[1807],M_list[1808],M_list[1809],M_list[1810],M_list[1811],M_list[1812],M_list[1813],M_list[1814],M_list[1815],M_list[1816],M_list[1817],M_list[1818],M_list[1819],M_list[1820],M_list[1821],M_list[1822],M_list[1823],M_list[1824],M_list[1825],M_list[1826],M_list[1827],M_list[1828],M_list[1829],M_list[1830],M_list[1831],M_list[1832],M_list[1833],M_list[1834],M_list[1835],M_list[1836],M_list[1837],M_list[1838],M_list[1839],M_list[1840],M_list[1841],M_list[1842],M_list[1843],M_list[1844],M_list[1845],M_list[1846],M_list[1847],M_list[1848],M_list[1849],M_list[1850],M_list[1851],M_list[1852],M_list[1853],M_list[1854],M_list[1855],M_list[1856],M_list[1857],M_list[1858],M_list[1859],M_list[1860],M_list[1861],M_list[1862],M_list[1863],M_list[1864],M_list[1865],M_list[1866],M_list[1867],M_list[1868],M_list[1869],M_list[1870],M_list[1871],M_list[1872],M_list[1873],M_list[1874],M_list[1875],M_list[1876],M_list[1877],M_list[1878],M_list[1879],M_list[1880],M_list[1881],M_list[1882],M_list[1883],M_list[1884],M_list[1885],M_list[1886],M_list[1887],M_list[1888],M_list[1889],M_list[1890],M_list[1891],M_list[1892],M_list[1893],M_list[1894],M_list[1895],M_list[1896],M_list[1897],M_list[1898],M_list[1899],M_list[1900],M_list[1901],M_list[1902],M_list[1903],M_list[1904],M_list[1905],M_list[1906],M_list[1907],M_list[1908],M_list[1909],M_list[1910],M_list[1911],M_list[1912],M_list[1913],M_list[1914],M_list[1915],M_list[1916],M_list[1917],M_list[1918],M_list[1919],M_list[1920],M_list[1921],M_list[1922],M_list[1923],M_list[1924],M_list[1925],M_list[1926],M_list[1927],M_list[1928],M_list[1929],M_list[1930],M_list[1931],M_list[1932],M_list[1933],M_list[1934],M_list[1935],M_list[1936],M_list[1937],M_list[1938],M_list[1939],M_list[1940],M_list[1941],M_list[1942],M_list[1943],M_list[1944],M_list[1945],M_list[1946],M_list[1947],M_list[1948],M_list[1949],M_list[1950],M_list[1951],M_list[1952],M_list[1953],M_list[1954],M_list[1955],M_list[1956],M_list[1957],M_list[1958],M_list[1959],M_list[1960],M_list[1961],M_list[1962],M_list[1963],M_list[1964],M_list[1965],M_list[1966],M_list[1967],M_list[1968],M_list[1969],M_list[1970],M_list[1971],M_list[1972],M_list[1973],M_list[1974],M_list[1975],M_list[1976],M_list[1977],M_list[1978],M_list[1979],M_list[1980],M_list[1981],M_list[1982],M_list[1983],M_list[1984],M_list[1985],M_list[1986],M_list[1987],M_list[1988],M_list[1989],M_list[1990],M_list[1991],M_list[1992],M_list[1993],M_list[1994],M_list[1995],M_list[1996],M_list[1997],M_list[1998],M_list[1999],M_list[2000],M_list[2001],M_list[2002],M_list[2003],M_list[2004],M_list[2005],M_list[2006],M_list[2007],M_list[2008],M_list[2009],M_list[2010],M_list[2011],M_list[2012],M_list[2013],M_list[2014],M_list[2015],M_list[2016],M_list[2017],M_list[2018],M_list[2019],M_list[2020],M_list[2021],M_list[2022],M_list[2023],M_list[2024],M_list[2025],M_list[2026],M_list[2027],M_list[2028],M_list[2029],M_list[2030],M_list[2031],M_list[2032],M_list[2033],M_list[2034],M_list[2035],M_list[2036],M_list[2037],M_list[2038],M_list[2039],M_list[2040],M_list[2041],M_list[2042],M_list[2043],M_list[2044],M_list[2045],M_list[2046],M_list[2047],M_list[2048],M_list[2049],M_list[2050],M_list[2051],M_list[2052],M_list[2053],M_list[2054],M_list[2055],M_list[2056],M_list[2057],M_list[2058],M_list[2059],M_list[2060],M_list[2061],M_list[2062],M_list[2063],M_list[2064],M_list[2065],M_list[2066],M_list[2067],M_list[2068],M_list[2069],M_list[2070],M_list[2071],M_list[2072],M_list[2073],M_list[2074],M_list[2075],M_list[2076],M_list[2077],M_list[2078],M_list[2079],M_list[2080],M_list[2081],M_list[2082],M_list[2083],M_list[2084],M_list[2085],M_list[2086],M_list[2087],M_list[2088],M_list[2089],M_list[2090],M_list[2091],M_list[2092],M_list[2093],M_list[2094],M_list[2095],M_list[2096],M_list[2097],M_list[2098],M_list[2099],M_list[2100],M_list[2101],M_list[2102],M_list[2103],M_list[2104],M_list[2105],M_list[2106],M_list[2107],M_list[2108],M_list[2109],M_list[2110],M_list[2111],M_list[2112],M_list[2113],M_list[2114],M_list[2115],M_list[2116],M_list[2117],M_list[2118],M_list[2119],M_list[2120],M_list[2121],M_list[2122],M_list[2123],M_list[2124],M_list[2125],M_list[2126],M_list[2127],M_list[2128],M_list[2129],M_list[2130],M_list[2131],M_list[2132],M_list[2133],M_list[2134],M_list[2135],M_list[2136],M_list[2137],M_list[2138],M_list[2139],M_list[2140],M_list[2141],M_list[2142],M_list[2143],M_list[2144],M_list[2145],M_list[2146],M_list[2147],M_list[2148],M_list[2149],M_list[2150],M_list[2151],M_list[2152],M_list[2153],M_list[2154],M_list[2155],M_list[2156],M_list[2157],M_list[2158],M_list[2159],M_list[2160],M_list[2161],M_list[2162],M_list[2163],M_list[2164],M_list[2165],M_list[2166],M_list[2167],M_list[2168],M_list[2169],M_list[2170],M_list[2171],M_list[2172],M_list[2173],M_list[2174],M_list[2175],M_list[2176],M_list[2177],M_list[2178],M_list[2179],M_list[2180],M_list[2181],M_list[2182],M_list[2183],M_list[2184],M_list[2185],M_list[2186],M_list[2187],M_list[2188],M_list[2189],M_list[2190],M_list[2191],M_list[2192],M_list[2193],M_list[2194],M_list[2195],M_list[2196],M_list[2197],M_list[2198],M_list[2199],M_list[2200],M_list[2201],M_list[2202],M_list[2203],M_list[2204],M_list[2205],M_list[2206],M_list[2207],M_list[2208],M_list[2209],M_list[2210],M_list[2211],M_list[2212],M_list[2213],M_list[2214],M_list[2215],M_list[2216],M_list[2217],M_list[2218],M_list[2219],M_list[2220],M_list[2221],M_list[2222],M_list[2223],M_list[2224],M_list[2225],M_list[2226],M_list[2227],M_list[2228],M_list[2229],M_list[2230],M_list[2231],M_list[2232],M_list[2233],M_list[2234],M_list[2235],M_list[2236],M_list[2237],M_list[2238],M_list[2239],M_list[2240],M_list[2241],M_list[2242],M_list[2243],M_list[2244],M_list[2245],M_list[2246],M_list[2247],M_list[2248],M_list[2249],M_list[2250],M_list[2251],M_list[2252],M_list[2253],M_list[2254],M_list[2255],M_list[2256],M_list[2257],M_list[2258],M_list[2259],M_list[2260],M_list[2261],M_list[2262],M_list[2263],M_list[2264],M_list[2265],M_list[2266],M_list[2267],M_list[2268],M_list[2269],M_list[2270],M_list[2271],M_list[2272],M_list[2273],M_list[2274],M_list[2275],M_list[2276],M_list[2277],M_list[2278],M_list[2279],M_list[2280],M_list[2281],M_list[2282],M_list[2283],M_list[2284],M_list[2285],M_list[2286],M_list[2287],M_list[2288],M_list[2289],M_list[2290],M_list[2291],M_list[2292],M_list[2293],M_list[2294],M_list[2295],M_list[2296],M_list[2297],M_list[2298],M_list[2299],M_list[2300],M_list[2301],M_list[2302],M_list[2303],M_list[2304],M_list[2305],M_list[2306],M_list[2307],M_list[2308],M_list[2309],M_list[2310],M_list[2311],M_list[2312],M_list[2313],M_list[2314],M_list[2315],M_list[2316],M_list[2317],M_list[2318],M_list[2319],M_list[2320],M_list[2321],M_list[2322],M_list[2323],M_list[2324],M_list[2325],M_list[2326],M_list[2327],M_list[2328],M_list[2329],M_list[2330],M_list[2331],M_list[2332],M_list[2333],M_list[2334],M_list[2335],M_list[2336],M_list[2337],M_list[2338],M_list[2339],M_list[2340],M_list[2341],M_list[2342],M_list[2343],M_list[2344],M_list[2345],M_list[2346],M_list[2347],M_list[2348],M_list[2349],M_list[2350],M_list[2351],M_list[2352],M_list[2353],M_list[2354],M_list[2355],M_list[2356],M_list[2357],M_list[2358],M_list[2359],M_list[2360],M_list[2361],M_list[2362],M_list[2363],M_list[2364],M_list[2365],M_list[2366],M_list[2367],M_list[2368],M_list[2369],M_list[2370],M_list[2371],M_list[2372],M_list[2373],M_list[2374],M_list[2375],M_list[2376],M_list[2377],M_list[2378],M_list[2379],M_list[2380],M_list[2381],M_list[2382],M_list[2383],M_list[2384],M_list[2385],M_list[2386],M_list[2387],M_list[2388],M_list[2389],M_list[2390],M_list[2391],M_list[2392],M_list[2393],M_list[2394],M_list[2395],M_list[2396],M_list[2397],M_list[2398],M_list[2399],M_list[2400],M_list[2401],M_list[2402],M_list[2403],M_list[2404],M_list[2405],M_list[2406],M_list[2407],M_list[2408],M_list[2409],M_list[2410],M_list[2411],M_list[2412],M_list[2413],M_list[2414],M_list[2415],M_list[2416],M_list[2417],M_list[2418],M_list[2419],M_list[2420],M_list[2421],M_list[2422],M_list[2423],M_list[2424],M_list[2425],M_list[2426],M_list[2427],M_list[2428],M_list[2429],M_list[2430],M_list[2431],M_list[2432],M_list[2433],M_list[2434],M_list[2435],M_list[2436],M_list[2437],M_list[2438],M_list[2439],M_list[2440],M_list[2441],M_list[2442],M_list[2443],M_list[2444],M_list[2445],M_list[2446],M_list[2447],M_list[2448],M_list[2449],M_list[2450],M_list[2451],M_list[2452],M_list[2453],M_list[2454],M_list[2455],M_list[2456],M_list[2457],M_list[2458],M_list[2459],M_list[2460],M_list[2461],M_list[2462],M_list[2463],M_list[2464],M_list[2465],M_list[2466],M_list[2467],M_list[2468],M_list[2469],M_list[2470],M_list[2471],M_list[2472],M_list[2473],M_list[2474],M_list[2475],M_list[2476],M_list[2477],M_list[2478],M_list[2479],M_list[2480],M_list[2481],M_list[2482],M_list[2483],M_list[2484],M_list[2485],M_list[2486],M_list[2487],M_list[2488],M_list[2489],M_list[2490],M_list[2491],M_list[2492],M_list[2493],M_list[2494],M_list[2495],M_list[2496],M_list[2497],M_list[2498],M_list[2499],M_list[2500],M_list[2501],M_list[2502],M_list[2503],M_list[2504],M_list[2505],M_list[2506],M_list[2507],M_list[2508],M_list[2509],M_list[2510],M_list[2511],M_list[2512],M_list[2513],M_list[2514],M_list[2515],M_list[2516],M_list[2517],M_list[2518],M_list[2519],M_list[2520],M_list[2521],M_list[2522],M_list[2523],M_list[2524],M_list[2525],M_list[2526],M_list[2527],M_list[2528],M_list[2529],M_list[2530],M_list[2531],M_list[2532],M_list[2533],M_list[2534],M_list[2535],M_list[2536],M_list[2537],M_list[2538],M_list[2539],M_list[2540],M_list[2541],M_list[2542],M_list[2543],M_list[2544],M_list[2545],M_list[2546],M_list[2547],M_list[2548],M_list[2549],M_list[2550],M_list[2551],M_list[2552],M_list[2553],M_list[2554],M_list[2555],M_list[2556],M_list[2557],M_list[2558],M_list[2559],M_list[2560],M_list[2561],M_list[2562],M_list[2563],M_list[2564],M_list[2565],M_list[2566],M_list[2567],M_list[2568],M_list[2569],M_list[2570],M_list[2571],M_list[2572],M_list[2573],M_list[2574],M_list[2575],M_list[2576],M_list[2577],M_list[2578],M_list[2579],M_list[2580],M_list[2581],M_list[2582],M_list[2583],M_list[2584],M_list[2585],M_list[2586],M_list[2587],M_list[2588],M_list[2589],M_list[2590],M_list[2591],M_list[2592],M_list[2593],M_list[2594],M_list[2595],M_list[2596],M_list[2597],M_list[2598],M_list[2599],M_list[2600],M_list[2601],M_list[2602],M_list[2603],M_list[2604],M_list[2605],M_list[2606],M_list[2607],M_list[2608],M_list[2609],M_list[2610],M_list[2611],M_list[2612],M_list[2613],M_list[2614],M_list[2615],M_list[2616],M_list[2617],M_list[2618],M_list[2619],M_list[2620],M_list[2621],M_list[2622],M_list[2623],M_list[2624],M_list[2625],M_list[2626],M_list[2627],M_list[2628],M_list[2629],M_list[2630],M_list[2631],M_list[2632],M_list[2633],M_list[2634],M_list[2635],M_list[2636],M_list[2637],M_list[2638],M_list[2639],M_list[2640],M_list[2641],M_list[2642],M_list[2643],M_list[2644],M_list[2645],M_list[2646],M_list[2647],M_list[2648],M_list[2649],M_list[2650],M_list[2651],M_list[2652],M_list[2653],M_list[2654],M_list[2655],M_list[2656],M_list[2657],M_list[2658],M_list[2659],M_list[2660],M_list[2661],M_list[2662],M_list[2663],M_list[2664],M_list[2665],M_list[2666],M_list[2667],M_list[2668],M_list[2669],M_list[2670],M_list[2671],M_list[2672],M_list[2673],M_list[2674],M_list[2675],M_list[2676],M_list[2677],M_list[2678],M_list[2679],M_list[2680],M_list[2681],M_list[2682],M_list[2683],M_list[2684],M_list[2685],M_list[2686],M_list[2687],M_list[2688],M_list[2689],M_list[2690],M_list[2691],M_list[2692],M_list[2693],M_list[2694],M_list[2695],M_list[2696],M_list[2697],M_list[2698],M_list[2699],M_list[2700],M_list[2701],M_list[2702],M_list[2703],M_list[2704],M_list[2705],M_list[2706],M_list[2707],M_list[2708],M_list[2709],M_list[2710],M_list[2711],M_list[2712],M_list[2713],M_list[2714],M_list[2715],M_list[2716],M_list[2717],M_list[2718],M_list[2719],M_list[2720],M_list[2721],M_list[2722],M_list[2723],M_list[2724],M_list[2725],M_list[2726],M_list[2727],M_list[2728],M_list[2729],M_list[2730],M_list[2731],M_list[2732],M_list[2733],M_list[2734],M_list[2735],M_list[2736],M_list[2737],M_list[2738],M_list[2739],M_list[2740],M_list[2741],M_list[2742],M_list[2743],M_list[2744],M_list[2745],M_list[2746],M_list[2747],M_list[2748],M_list[2749],M_list[2750],M_list[2751],M_list[2752],M_list[2753],M_list[2754],M_list[2755],M_list[2756],M_list[2757],M_list[2758],M_list[2759],M_list[2760],M_list[2761],M_list[2762],M_list[2763],M_list[2764],M_list[2765],M_list[2766],M_list[2767],M_list[2768],M_list[2769],M_list[2770],M_list[2771],M_list[2772],M_list[2773],M_list[2774],M_list[2775],M_list[2776],M_list[2777],M_list[2778],M_list[2779],M_list[2780],M_list[2781],M_list[2782],M_list[2783],M_list[2784],M_list[2785],M_list[2786],M_list[2787],M_list[2788],M_list[2789],M_list[2790],M_list[2791],M_list[2792],M_list[2793],M_list[2794],M_list[2795],M_list[2796],M_list[2797],M_list[2798],M_list[2799],M_list[2800],M_list[2801],M_list[2802],M_list[2803],M_list[2804],M_list[2805],M_list[2806],M_list[2807],M_list[2808],M_list[2809],M_list[2810],M_list[2811],M_list[2812],M_list[2813],M_list[2814],M_list[2815],M_list[2816],M_list[2817],M_list[2818],M_list[2819],M_list[2820],M_list[2821],M_list[2822],M_list[2823],M_list[2824],M_list[2825],M_list[2826],M_list[2827],M_list[2828],M_list[2829],M_list[2830],M_list[2831],M_list[2832],M_list[2833],M_list[2834],M_list[2835],M_list[2836],M_list[2837],M_list[2838],M_list[2839],M_list[2840],M_list[2841],M_list[2842],M_list[2843],M_list[2844],M_list[2845],M_list[2846],M_list[2847],M_list[2848],M_list[2849],M_list[2850],M_list[2851],M_list[2852],M_list[2853],M_list[2854],M_list[2855],M_list[2856],M_list[2857],M_list[2858],M_list[2859],M_list[2860],M_list[2861],M_list[2862],M_list[2863],M_list[2864],M_list[2865],M_list[2866],M_list[2867],M_list[2868],M_list[2869],M_list[2870],M_list[2871],M_list[2872],M_list[2873],M_list[2874],M_list[2875],M_list[2876],M_list[2877],M_list[2878],M_list[2879],M_list[2880],M_list[2881],M_list[2882],M_list[2883],M_list[2884],M_list[2885],M_list[2886],M_list[2887],M_list[2888],M_list[2889],M_list[2890],M_list[2891],M_list[2892],M_list[2893],M_list[2894],M_list[2895],M_list[2896],M_list[2897],M_list[2898],M_list[2899],M_list[2900],M_list[2901],M_list[2902],M_list[2903],M_list[2904],M_list[2905],M_list[2906],M_list[2907],M_list[2908],M_list[2909],M_list[2910],M_list[2911],M_list[2912],M_list[2913],M_list[2914],M_list[2915],M_list[2916],M_list[2917],M_list[2918],M_list[2919],M_list[2920],M_list[2921],M_list[2922],M_list[2923],M_list[2924],M_list[2925],M_list[2926],M_list[2927],M_list[2928],M_list[2929],M_list[2930],M_list[2931],M_list[2932],M_list[2933],M_list[2934],M_list[2935],M_list[2936],M_list[2937],M_list[2938],M_list[2939],M_list[2940],M_list[2941],M_list[2942],M_list[2943],M_list[2944],M_list[2945],M_list[2946],M_list[2947],M_list[2948],M_list[2949],M_list[2950],M_list[2951],M_list[2952],M_list[2953],M_list[2954],M_list[2955],M_list[2956],M_list[2957],M_list[2958],M_list[2959],M_list[2960],M_list[2961],M_list[2962],M_list[2963],M_list[2964],M_list[2965],M_list[2966],M_list[2967],M_list[2968],M_list[2969],M_list[2970],M_list[2971],M_list[2972],M_list[2973],M_list[2974],M_list[2975],M_list[2976],M_list[2977],M_list[2978],M_list[2979],M_list[2980],M_list[2981],M_list[2982],M_list[2983],M_list[2984],M_list[2985],M_list[2986],M_list[2987],M_list[2988],M_list[2989],M_list[2990],M_list[2991],M_list[2992],M_list[2993],M_list[2994],M_list[2995],M_list[2996],M_list[2997],M_list[2998],M_list[2999],M_list[3000],M_list[3001],M_list[3002],M_list[3003],M_list[3004],M_list[3005],M_list[3006],M_list[3007],M_list[3008],M_list[3009],M_list[3010],M_list[3011],M_list[3012],M_list[3013],M_list[3014],M_list[3015],M_list[3016],M_list[3017],M_list[3018],M_list[3019],M_list[3020],M_list[3021],M_list[3022],M_list[3023],M_list[3024],M_list[3025],M_list[3026],M_list[3027],M_list[3028],M_list[3029],M_list[3030],M_list[3031],M_list[3032],M_list[3033],M_list[3034],M_list[3035],M_list[3036],M_list[3037],M_list[3038],M_list[3039],M_list[3040],M_list[3041],M_list[3042],M_list[3043],M_list[3044],M_list[3045],M_list[3046],M_list[3047],M_list[3048],M_list[3049],M_list[3050],M_list[3051],M_list[3052],M_list[3053],M_list[3054],M_list[3055],M_list[3056],M_list[3057],M_list[3058],M_list[3059],M_list[3060],M_list[3061],M_list[3062],M_list[3063],M_list[3064],M_list[3065],M_list[3066],M_list[3067],M_list[3068],M_list[3069],M_list[3070],M_list[3071],M_list[3072],M_list[3073],M_list[3074],M_list[3075],M_list[3076],M_list[3077],M_list[3078],M_list[3079],M_list[3080],M_list[3081],M_list[3082],M_list[3083],M_list[3084],M_list[3085],M_list[3086],M_list[3087],M_list[3088],M_list[3089],M_list[3090],M_list[3091],M_list[3092],M_list[3093],M_list[3094],M_list[3095],M_list[3096],M_list[3097],M_list[3098],M_list[3099],M_list[3100],M_list[3101],M_list[3102],M_list[3103],M_list[3104],M_list[3105],M_list[3106],M_list[3107],M_list[3108],M_list[3109],M_list[3110],M_list[3111],M_list[3112],M_list[3113],M_list[3114],M_list[3115],M_list[3116],M_list[3117],M_list[3118],M_list[3119],M_list[3120],M_list[3121],M_list[3122],M_list[3123],M_list[3124],M_list[3125],M_list[3126],M_list[3127],M_list[3128],M_list[3129],M_list[3130],M_list[3131],M_list[3132],M_list[3133],M_list[3134],M_list[3135],M_list[3136],M_list[3137],M_list[3138],M_list[3139],M_list[3140],M_list[3141],M_list[3142],M_list[3143],M_list[3144],M_list[3145],M_list[3146],M_list[3147],M_list[3148],M_list[3149],M_list[3150],M_list[3151],M_list[3152],M_list[3153],M_list[3154],M_list[3155],M_list[3156],M_list[3157],M_list[3158],M_list[3159],M_list[3160],M_list[3161],M_list[3162],M_list[3163],M_list[3164],M_list[3165],M_list[3166],M_list[3167],M_list[3168],M_list[3169],M_list[3170],M_list[3171],M_list[3172],M_list[3173],M_list[3174],M_list[3175],M_list[3176],M_list[3177],M_list[3178],M_list[3179],M_list[3180],M_list[3181],M_list[3182],M_list[3183],M_list[3184],M_list[3185],M_list[3186],M_list[3187],M_list[3188],M_list[3189],M_list[3190],M_list[3191],M_list[3192],M_list[3193],M_list[3194],M_list[3195],M_list[3196],M_list[3197],M_list[3198],M_list[3199],M_list[3200],M_list[3201],M_list[3202],M_list[3203],M_list[3204],M_list[3205],M_list[3206],M_list[3207],M_list[3208],M_list[3209],M_list[3210],M_list[3211],M_list[3212],M_list[3213],M_list[3214],M_list[3215],M_list[3216],M_list[3217],M_list[3218],M_list[3219],M_list[3220],M_list[3221],M_list[3222],M_list[3223],M_list[3224],M_list[3225],M_list[3226],M_list[3227],M_list[3228],M_list[3229],M_list[3230],M_list[3231],M_list[3232],M_list[3233],M_list[3234],M_list[3235],M_list[3236],M_list[3237],M_list[3238],M_list[3239],M_list[3240],M_list[3241],M_list[3242],M_list[3243],M_list[3244],M_list[3245],M_list[3246],M_list[3247],M_list[3248],M_list[3249],M_list[3250],M_list[3251],M_list[3252],M_list[3253],M_list[3254],M_list[3255],M_list[3256],M_list[3257],M_list[3258],M_list[3259],M_list[3260],M_list[3261],M_list[3262],M_list[3263],M_list[3264],M_list[3265],M_list[3266],M_list[3267],M_list[3268],M_list[3269],M_list[3270],M_list[3271],M_list[3272],M_list[3273],M_list[3274],M_list[3275],M_list[3276],M_list[3277],M_list[3278],M_list[3279],M_list[3280],M_list[3281],M_list[3282],M_list[3283],M_list[3284],M_list[3285],M_list[3286],M_list[3287],M_list[3288],M_list[3289],M_list[3290],M_list[3291],M_list[3292],M_list[3293],M_list[3294],M_list[3295],M_list[3296],M_list[3297],M_list[3298],M_list[3299],M_list[3300],M_list[3301],M_list[3302],M_list[3303],M_list[3304],M_list[3305],M_list[3306],M_list[3307],M_list[3308],M_list[3309],M_list[3310],M_list[3311],M_list[3312],M_list[3313],M_list[3314],M_list[3315],M_list[3316],M_list[3317],M_list[3318],M_list[3319],M_list[3320],M_list[3321],M_list[3322],M_list[3323],M_list[3324],M_list[3325],M_list[3326],M_list[3327],M_list[3328],M_list[3329],M_list[3330],M_list[3331],M_list[3332],M_list[3333],M_list[3334],M_list[3335],M_list[3336],M_list[3337],M_list[3338],M_list[3339],M_list[3340],M_list[3341],M_list[3342],M_list[3343],M_list[3344],M_list[3345],M_list[3346],M_list[3347],M_list[3348],M_list[3349],M_list[3350],M_list[3351],M_list[3352],M_list[3353],M_list[3354],M_list[3355],M_list[3356],M_list[3357],M_list[3358],M_list[3359],M_list[3360],M_list[3361],M_list[3362],M_list[3363],M_list[3364],M_list[3365],M_list[3366],M_list[3367],M_list[3368],M_list[3369],M_list[3370],M_list[3371],M_list[3372],M_list[3373],M_list[3374],M_list[3375],M_list[3376],M_list[3377],M_list[3378],M_list[3379],M_list[3380],M_list[3381],M_list[3382],M_list[3383],M_list[3384],M_list[3385],M_list[3386],M_list[3387],M_list[3388],M_list[3389],M_list[3390],M_list[3391],M_list[3392],M_list[3393],M_list[3394],M_list[3395],M_list[3396],M_list[3397],M_list[3398],M_list[3399],M_list[3400],M_list[3401],M_list[3402],M_list[3403],M_list[3404],M_list[3405],M_list[3406],M_list[3407],M_list[3408],M_list[3409],M_list[3410],M_list[3411],M_list[3412],M_list[3413],M_list[3414],M_list[3415],M_list[3416],M_list[3417],M_list[3418],M_list[3419],M_list[3420],M_list[3421],M_list[3422],M_list[3423],M_list[3424],M_list[3425],M_list[3426],M_list[3427],M_list[3428],M_list[3429],M_list[3430],M_list[3431],M_list[3432],M_list[3433],M_list[3434],M_list[3435],M_list[3436],M_list[3437],M_list[3438],M_list[3439],M_list[3440],M_list[3441],M_list[3442],M_list[3443],M_list[3444],M_list[3445],M_list[3446],M_list[3447],M_list[3448],M_list[3449],M_list[3450],M_list[3451],M_list[3452],M_list[3453],M_list[3454],M_list[3455],M_list[3456],M_list[3457],M_list[3458],M_list[3459],M_list[3460],M_list[3461],M_list[3462],M_list[3463],M_list[3464],M_list[3465],M_list[3466],M_list[3467],M_list[3468],M_list[3469],M_list[3470],M_list[3471],M_list[3472],M_list[3473],M_list[3474],M_list[3475],M_list[3476],M_list[3477],M_list[3478],M_list[3479],M_list[3480],M_list[3481],M_list[3482],M_list[3483],M_list[3484],M_list[3485],M_list[3486],M_list[3487],M_list[3488],M_list[3489],M_list[3490],M_list[3491],M_list[3492],M_list[3493],M_list[3494],M_list[3495],M_list[3496],M_list[3497],M_list[3498],M_list[3499],M_list[3500],M_list[3501],M_list[3502],M_list[3503],M_list[3504],M_list[3505],M_list[3506],M_list[3507],M_list[3508],M_list[3509],M_list[3510],M_list[3511],M_list[3512],M_list[3513],M_list[3514],M_list[3515],M_list[3516],M_list[3517],M_list[3518],M_list[3519],M_list[3520],M_list[3521],M_list[3522],M_list[3523],M_list[3524],M_list[3525],M_list[3526],M_list[3527],M_list[3528],M_list[3529],M_list[3530],M_list[3531],M_list[3532],M_list[3533],M_list[3534],M_list[3535],M_list[3536],M_list[3537],M_list[3538],M_list[3539],M_list[3540],M_list[3541],M_list[3542],M_list[3543],M_list[3544],M_list[3545],M_list[3546],M_list[3547],M_list[3548],M_list[3549],M_list[3550],M_list[3551],M_list[3552],M_list[3553],M_list[3554],M_list[3555],M_list[3556],M_list[3557],M_list[3558],M_list[3559],M_list[3560],M_list[3561],M_list[3562],M_list[3563],M_list[3564],M_list[3565],M_list[3566],M_list[3567],M_list[3568],M_list[3569],M_list[3570],M_list[3571],M_list[3572],M_list[3573],M_list[3574],M_list[3575],M_list[3576],M_list[3577],M_list[3578],M_list[3579],M_list[3580],M_list[3581],M_list[3582],M_list[3583],M_list[3584],M_list[3585],M_list[3586],M_list[3587],M_list[3588],M_list[3589],M_list[3590],M_list[3591],M_list[3592],M_list[3593],M_list[3594],M_list[3595],M_list[3596],M_list[3597],M_list[3598],M_list[3599],M_list[3600],M_list[3601],M_list[3602],M_list[3603],M_list[3604],M_list[3605],M_list[3606],M_list[3607],M_list[3608],M_list[3609],M_list[3610],M_list[3611],M_list[3612],M_list[3613],M_list[3614],M_list[3615],M_list[3616],M_list[3617],M_list[3618],M_list[3619],M_list[3620],M_list[3621],M_list[3622],M_list[3623],M_list[3624],M_list[3625],M_list[3626],M_list[3627],M_list[3628],M_list[3629],M_list[3630],M_list[3631],M_list[3632],M_list[3633],M_list[3634],M_list[3635],M_list[3636],M_list[3637],M_list[3638],M_list[3639],M_list[3640],M_list[3641],M_list[3642],M_list[3643],M_list[3644],M_list[3645],M_list[3646],M_list[3647],M_list[3648],M_list[3649],M_list[3650],M_list[3651],M_list[3652],M_list[3653],M_list[3654],M_list[3655],M_list[3656],M_list[3657],M_list[3658],M_list[3659],M_list[3660],M_list[3661],M_list[3662],M_list[3663],M_list[3664],M_list[3665],M_list[3666],M_list[3667],M_list[3668],M_list[3669],M_list[3670],M_list[3671],M_list[3672],M_list[3673],M_list[3674],M_list[3675],M_list[3676],M_list[3677],M_list[3678],M_list[3679],M_list[3680],M_list[3681],M_list[3682],M_list[3683],M_list[3684],M_list[3685],M_list[3686],M_list[3687],M_list[3688],M_list[3689],M_list[3690],M_list[3691],M_list[3692],M_list[3693],M_list[3694],M_list[3695],M_list[3696],M_list[3697],M_list[3698],M_list[3699],M_list[3700],M_list[3701],M_list[3702],M_list[3703],M_list[3704],M_list[3705],M_list[3706],M_list[3707],M_list[3708],M_list[3709],M_list[3710],M_list[3711],M_list[3712],M_list[3713],M_list[3714],M_list[3715],M_list[3716],M_list[3717],M_list[3718],M_list[3719],M_list[3720],M_list[3721],M_list[3722],M_list[3723],M_list[3724],M_list[3725],M_list[3726],M_list[3727],M_list[3728],M_list[3729],M_list[3730],M_list[3731],M_list[3732],M_list[3733],M_list[3734],M_list[3735],M_list[3736],M_list[3737],M_list[3738],M_list[3739],M_list[3740],M_list[3741],M_list[3742],M_list[3743],M_list[3744],M_list[3745],M_list[3746],M_list[3747],M_list[3748],M_list[3749],M_list[3750],M_list[3751],M_list[3752],M_list[3753],M_list[3754],M_list[3755],M_list[3756],M_list[3757],M_list[3758],M_list[3759],M_list[3760],M_list[3761],M_list[3762],M_list[3763],M_list[3764],M_list[3765],M_list[3766],M_list[3767],M_list[3768],M_list[3769],M_list[3770],M_list[3771],M_list[3772],M_list[3773],M_list[3774],M_list[3775],M_list[3776],M_list[3777],M_list[3778],M_list[3779],M_list[3780],M_list[3781],M_list[3782],M_list[3783],M_list[3784],M_list[3785],M_list[3786],M_list[3787],M_list[3788],M_list[3789],M_list[3790],M_list[3791],M_list[3792],M_list[3793],M_list[3794],M_list[3795],M_list[3796],M_list[3797],M_list[3798],M_list[3799],M_list[3800],M_list[3801],M_list[3802],M_list[3803],M_list[3804],M_list[3805],M_list[3806],M_list[3807],M_list[3808],M_list[3809],M_list[3810],M_list[3811],M_list[3812],M_list[3813],M_list[3814],M_list[3815],M_list[3816],M_list[3817],M_list[3818],M_list[3819],M_list[3820],M_list[3821],M_list[3822],M_list[3823],M_list[3824],M_list[3825],M_list[3826],M_list[3827],M_list[3828],M_list[3829],M_list[3830],M_list[3831],M_list[3832],M_list[3833],M_list[3834],M_list[3835],M_list[3836],M_list[3837],M_list[3838],M_list[3839],M_list[3840],M_list[3841],M_list[3842],M_list[3843],M_list[3844],M_list[3845],M_list[3846],M_list[3847],M_list[3848],M_list[3849],M_list[3850],M_list[3851],M_list[3852],M_list[3853],M_list[3854],M_list[3855],M_list[3856],M_list[3857],M_list[3858],M_list[3859],M_list[3860],M_list[3861],M_list[3862],M_list[3863],M_list[3864],M_list[3865],M_list[3866],M_list[3867],M_list[3868],M_list[3869],M_list[3870],M_list[3871],M_list[3872],M_list[3873],M_list[3874],M_list[3875],M_list[3876],M_list[3877],M_list[3878],M_list[3879],M_list[3880],M_list[3881],M_list[3882],M_list[3883],M_list[3884],M_list[3885],M_list[3886],M_list[3887],M_list[3888],M_list[3889],M_list[3890],M_list[3891],M_list[3892],M_list[3893],M_list[3894],M_list[3895],M_list[3896],M_list[3897],M_list[3898],M_list[3899],M_list[3900],M_list[3901],M_list[3902],M_list[3903],M_list[3904],M_list[3905],M_list[3906],M_list[3907],M_list[3908],M_list[3909],M_list[3910],M_list[3911],M_list[3912],M_list[3913],M_list[3914],M_list[3915],M_list[3916],M_list[3917],M_list[3918],M_list[3919],M_list[3920],M_list[3921],M_list[3922],M_list[3923],M_list[3924],M_list[3925],M_list[3926],M_list[3927],M_list[3928],M_list[3929],M_list[3930],M_list[3931],M_list[3932],M_list[3933],M_list[3934],M_list[3935],M_list[3936],M_list[3937],M_list[3938],M_list[3939],M_list[3940],M_list[3941],M_list[3942],M_list[3943],M_list[3944],M_list[3945],M_list[3946],M_list[3947],M_list[3948],M_list[3949],M_list[3950],M_list[3951],M_list[3952],M_list[3953],M_list[3954],M_list[3955],M_list[3956],M_list[3957],M_list[3958],M_list[3959],M_list[3960],M_list[3961],M_list[3962],M_list[3963],M_list[3964],M_list[3965],M_list[3966],M_list[3967],M_list[3968],M_list[3969],M_list[3970],M_list[3971],M_list[3972],M_list[3973],M_list[3974],M_list[3975],M_list[3976],M_list[3977],M_list[3978],M_list[3979],M_list[3980],M_list[3981],M_list[3982],M_list[3983],M_list[3984],M_list[3985],M_list[3986],M_list[3987],M_list[3988],M_list[3989],M_list[3990],M_list[3991],M_list[3992],M_list[3993],M_list[3994],M_list[3995],M_list[3996],M_list[3997],M_list[3998],M_list[3999],M_list[4000],M_list[4001],M_list[4002],M_list[4003],M_list[4004],M_list[4005],M_list[4006],M_list[4007],M_list[4008],M_list[4009],M_list[4010],M_list[4011],M_list[4012],M_list[4013],M_list[4014],M_list[4015],M_list[4016],M_list[4017],M_list[4018],M_list[4019],M_list[4020],M_list[4021],M_list[4022],M_list[4023],M_list[4024],M_list[4025],M_list[4026],M_list[4027],M_list[4028],M_list[4029],M_list[4030],M_list[4031],M_list[4032],M_list[4033],M_list[4034],M_list[4035],M_list[4036],M_list[4037],M_list[4038],M_list[4039],M_list[4040],M_list[4041],M_list[4042],M_list[4043],M_list[4044],M_list[4045],M_list[4046],M_list[4047],M_list[4048],M_list[4049],M_list[4050],M_list[4051],M_list[4052],M_list[4053],M_list[4054],M_list[4055],M_list[4056],M_list[4057],M_list[4058],M_list[4059],M_list[4060],M_list[4061],M_list[4062],M_list[4063],M_list[4064],M_list[4065],M_list[4066],M_list[4067],M_list[4068],M_list[4069],M_list[4070],M_list[4071],M_list[4072],M_list[4073],M_list[4074],M_list[4075],M_list[4076],M_list[4077],M_list[4078],M_list[4079],M_list[4080],M_list[4081],M_list[4082],M_list[4083],M_list[4084],M_list[4085],M_list[4086],M_list[4087],M_list[4088],M_list[4089],M_list[4090],M_list[4091],M_list[4092],M_list[4093],M_list[4094],M_list[4095],M_list[4096],M_list[4097],M_list[4098],M_list[4099],M_list[4100],M_list[4101],M_list[4102],M_list[4103],M_list[4104],M_list[4105],M_list[4106],M_list[4107],M_list[4108],M_list[4109],M_list[4110],M_list[4111],M_list[4112],M_list[4113],M_list[4114],M_list[4115],M_list[4116],M_list[4117],M_list[4118],M_list[4119],M_list[4120],M_list[4121],M_list[4122],M_list[4123],M_list[4124],M_list[4125],M_list[4126],M_list[4127],M_list[4128],M_list[4129],M_list[4130],M_list[4131],M_list[4132],M_list[4133],M_list[4134],M_list[4135],M_list[4136],M_list[4137],M_list[4138],M_list[4139],M_list[4140],M_list[4141],M_list[4142],M_list[4143],M_list[4144],M_list[4145],M_list[4146],M_list[4147],M_list[4148],M_list[4149],M_list[4150],M_list[4151],M_list[4152],M_list[4153],M_list[4154],M_list[4155],M_list[4156],M_list[4157],M_list[4158],M_list[4159],M_list[4160],M_list[4161],M_list[4162],M_list[4163],M_list[4164],M_list[4165],M_list[4166],M_list[4167],M_list[4168],M_list[4169],M_list[4170],M_list[4171],M_list[4172],M_list[4173],M_list[4174],M_list[4175],M_list[4176],M_list[4177],M_list[4178],M_list[4179],M_list[4180],M_list[4181],M_list[4182],M_list[4183],M_list[4184],M_list[4185],M_list[4186],M_list[4187],M_list[4188],M_list[4189],M_list[4190],M_list[4191],M_list[4192],M_list[4193],M_list[4194],M_list[4195],M_list[4196],M_list[4197],M_list[4198],M_list[4199],M_list[4200],M_list[4201],M_list[4202],M_list[4203],M_list[4204],M_list[4205],M_list[4206],M_list[4207],M_list[4208],M_list[4209],M_list[4210],M_list[4211],M_list[4212],M_list[4213],M_list[4214],M_list[4215],M_list[4216],M_list[4217],M_list[4218],M_list[4219],M_list[4220],M_list[4221],M_list[4222],M_list[4223],M_list[4224],M_list[4225],M_list[4226],M_list[4227],M_list[4228],M_list[4229],M_list[4230],M_list[4231],M_list[4232],M_list[4233],M_list[4234],M_list[4235],M_list[4236],M_list[4237],M_list[4238],M_list[4239],M_list[4240],M_list[4241],M_list[4242],M_list[4243],M_list[4244],M_list[4245],M_list[4246],M_list[4247],M_list[4248],M_list[4249],M_list[4250],M_list[4251],M_list[4252],M_list[4253],M_list[4254],M_list[4255],M_list[4256],M_list[4257],M_list[4258],M_list[4259],M_list[4260],M_list[4261],M_list[4262],M_list[4263],M_list[4264],M_list[4265],M_list[4266],M_list[4267],M_list[4268],M_list[4269],M_list[4270],M_list[4271],M_list[4272],M_list[4273],M_list[4274],M_list[4275],M_list[4276],M_list[4277],M_list[4278],M_list[4279],M_list[4280],M_list[4281],M_list[4282],M_list[4283],M_list[4284],M_list[4285],M_list[4286],M_list[4287],M_list[4288],M_list[4289],M_list[4290],M_list[4291],M_list[4292],M_list[4293],M_list[4294],M_list[4295],M_list[4296],M_list[4297],M_list[4298],M_list[4299],M_list[4300],M_list[4301],M_list[4302],M_list[4303],M_list[4304],M_list[4305],M_list[4306],M_list[4307],M_list[4308],M_list[4309],M_list[4310],M_list[4311],M_list[4312],M_list[4313],M_list[4314],M_list[4315],M_list[4316],M_list[4317],M_list[4318],M_list[4319],M_list[4320],M_list[4321],M_list[4322],M_list[4323],M_list[4324],M_list[4325],M_list[4326],M_list[4327],M_list[4328],M_list[4329],M_list[4330],M_list[4331],M_list[4332],M_list[4333],M_list[4334],M_list[4335],M_list[4336],M_list[4337],M_list[4338],M_list[4339],M_list[4340],M_list[4341],M_list[4342],M_list[4343],M_list[4344],M_list[4345],M_list[4346],M_list[4347],M_list[4348],M_list[4349],M_list[4350],M_list[4351],M_list[4352],M_list[4353],M_list[4354],M_list[4355],M_list[4356],M_list[4357],M_list[4358],M_list[4359],M_list[4360],M_list[4361],M_list[4362],M_list[4363],M_list[4364],M_list[4365],M_list[4366],M_list[4367],M_list[4368],M_list[4369],M_list[4370],M_list[4371],M_list[4372],M_list[4373],M_list[4374],M_list[4375],M_list[4376],M_list[4377],M_list[4378],M_list[4379],M_list[4380],M_list[4381],M_list[4382],M_list[4383],M_list[4384],M_list[4385],M_list[4386],M_list[4387],M_list[4388],M_list[4389],M_list[4390],M_list[4391],M_list[4392],M_list[4393],M_list[4394],M_list[4395],M_list[4396],M_list[4397],M_list[4398],M_list[4399],M_list[4400],M_list[4401],M_list[4402],M_list[4403],M_list[4404],M_list[4405],M_list[4406],M_list[4407],M_list[4408],M_list[4409],M_list[4410],M_list[4411],M_list[4412],M_list[4413],M_list[4414],M_list[4415],M_list[4416],M_list[4417],M_list[4418],M_list[4419],M_list[4420],M_list[4421],M_list[4422],M_list[4423],M_list[4424],M_list[4425],M_list[4426],M_list[4427],M_list[4428],M_list[4429],M_list[4430],M_list[4431],M_list[4432],M_list[4433],M_list[4434],M_list[4435],M_list[4436],M_list[4437],M_list[4438],M_list[4439],M_list[4440],M_list[4441],M_list[4442],M_list[4443],M_list[4444],M_list[4445],M_list[4446],M_list[4447],M_list[4448],M_list[4449],M_list[4450],M_list[4451],M_list[4452],M_list[4453],M_list[4454],M_list[4455],M_list[4456],M_list[4457],M_list[4458],M_list[4459],M_list[4460],M_list[4461],M_list[4462],M_list[4463],M_list[4464],M_list[4465],M_list[4466],M_list[4467],M_list[4468],M_list[4469],M_list[4470],M_list[4471],M_list[4472],M_list[4473],M_list[4474],M_list[4475],M_list[4476],M_list[4477],M_list[4478],M_list[4479],M_list[4480],M_list[4481],M_list[4482],M_list[4483],M_list[4484],M_list[4485],M_list[4486],M_list[4487],M_list[4488],M_list[4489],M_list[4490],M_list[4491],M_list[4492],M_list[4493],M_list[4494],M_list[4495],M_list[4496],M_list[4497],M_list[4498],M_list[4499],M_list[4500],M_list[4501],M_list[4502],M_list[4503],M_list[4504],M_list[4505],M_list[4506],M_list[4507],M_list[4508],M_list[4509],M_list[4510],M_list[4511],M_list[4512],M_list[4513],M_list[4514],M_list[4515],M_list[4516],M_list[4517],M_list[4518],M_list[4519],M_list[4520],M_list[4521],M_list[4522],M_list[4523],M_list[4524],M_list[4525],M_list[4526],M_list[4527],M_list[4528],M_list[4529],M_list[4530],M_list[4531],M_list[4532],M_list[4533],M_list[4534],M_list[4535],M_list[4536],M_list[4537],M_list[4538],M_list[4539],M_list[4540],M_list[4541],M_list[4542],M_list[4543],M_list[4544],M_list[4545],M_list[4546],M_list[4547],M_list[4548],M_list[4549],M_list[4550],M_list[4551],M_list[4552],M_list[4553],M_list[4554],M_list[4555],M_list[4556],M_list[4557],M_list[4558],M_list[4559],M_list[4560],M_list[4561],M_list[4562],M_list[4563],M_list[4564],M_list[4565],M_list[4566],M_list[4567],M_list[4568],M_list[4569],M_list[4570],M_list[4571],M_list[4572],M_list[4573],M_list[4574],M_list[4575],M_list[4576],M_list[4577],M_list[4578],M_list[4579],M_list[4580],M_list[4581],M_list[4582],M_list[4583],M_list[4584],M_list[4585],M_list[4586],M_list[4587],M_list[4588],M_list[4589],M_list[4590],M_list[4591],M_list[4592],M_list[4593],M_list[4594],M_list[4595],M_list[4596],M_list[4597],M_list[4598],M_list[4599],M_list[4600],M_list[4601],M_list[4602],M_list[4603],M_list[4604],M_list[4605],M_list[4606],M_list[4607],M_list[4608],M_list[4609],M_list[4610],M_list[4611],M_list[4612],M_list[4613],M_list[4614],M_list[4615],M_list[4616],M_list[4617],M_list[4618],M_list[4619],M_list[4620],M_list[4621],M_list[4622],M_list[4623],M_list[4624],M_list[4625],M_list[4626],M_list[4627],M_list[4628],M_list[4629],M_list[4630],M_list[4631],M_list[4632],M_list[4633],M_list[4634],M_list[4635],M_list[4636],M_list[4637],M_list[4638],M_list[4639],M_list[4640],M_list[4641],M_list[4642],M_list[4643],M_list[4644],M_list[4645],M_list[4646],M_list[4647],M_list[4648],M_list[4649],M_list[4650],M_list[4651],M_list[4652],M_list[4653],M_list[4654],M_list[4655],M_list[4656],M_list[4657],M_list[4658],M_list[4659],M_list[4660],M_list[4661],M_list[4662],M_list[4663],M_list[4664],M_list[4665],M_list[4666],M_list[4667],M_list[4668],M_list[4669],M_list[4670],M_list[4671],M_list[4672],M_list[4673],M_list[4674],M_list[4675],M_list[4676],M_list[4677],M_list[4678],M_list[4679],M_list[4680],M_list[4681],M_list[4682],M_list[4683],M_list[4684],M_list[4685],M_list[4686],M_list[4687],M_list[4688],M_list[4689],M_list[4690],M_list[4691],M_list[4692],M_list[4693],M_list[4694],M_list[4695],M_list[4696],M_list[4697],M_list[4698],M_list[4699],M_list[4700],M_list[4701],M_list[4702],M_list[4703],M_list[4704],M_list[4705],M_list[4706],M_list[4707],M_list[4708],M_list[4709],M_list[4710],M_list[4711],M_list[4712],M_list[4713],M_list[4714],M_list[4715],M_list[4716],M_list[4717],M_list[4718],M_list[4719],M_list[4720],M_list[4721],M_list[4722],M_list[4723],M_list[4724],M_list[4725],M_list[4726],M_list[4727],M_list[4728],M_list[4729],M_list[4730],M_list[4731],M_list[4732],M_list[4733],M_list[4734],M_list[4735],M_list[4736],M_list[4737],M_list[4738],M_list[4739],M_list[4740],M_list[4741],M_list[4742],M_list[4743],M_list[4744],M_list[4745],M_list[4746],M_list[4747],M_list[4748],M_list[4749],M_list[4750],M_list[4751],M_list[4752],M_list[4753],M_list[4754],M_list[4755],M_list[4756],M_list[4757],M_list[4758],M_list[4759],M_list[4760],M_list[4761],M_list[4762],M_list[4763],M_list[4764],M_list[4765],M_list[4766],M_list[4767],M_list[4768],M_list[4769],M_list[4770],M_list[4771],M_list[4772],M_list[4773],M_list[4774],M_list[4775],M_list[4776],M_list[4777],M_list[4778],M_list[4779],M_list[4780],M_list[4781],M_list[4782],M_list[4783],M_list[4784],M_list[4785],M_list[4786],M_list[4787],M_list[4788],M_list[4789],M_list[4790],M_list[4791],M_list[4792],M_list[4793],M_list[4794],M_list[4795],M_list[4796],M_list[4797],M_list[4798],M_list[4799],M_list[4800],M_list[4801],M_list[4802],M_list[4803],M_list[4804],M_list[4805],M_list[4806],M_list[4807],M_list[4808],M_list[4809],M_list[4810],M_list[4811],M_list[4812],M_list[4813],M_list[4814],M_list[4815],M_list[4816],M_list[4817],M_list[4818],M_list[4819],M_list[4820],M_list[4821],M_list[4822],M_list[4823],M_list[4824],M_list[4825],M_list[4826],M_list[4827],M_list[4828],M_list[4829],M_list[4830],M_list[4831],M_list[4832],M_list[4833],M_list[4834],M_list[4835],M_list[4836],M_list[4837],M_list[4838],M_list[4839],M_list[4840],M_list[4841],M_list[4842],M_list[4843],M_list[4844],M_list[4845],M_list[4846],M_list[4847],M_list[4848],M_list[4849],M_list[4850],M_list[4851],M_list[4852],M_list[4853],M_list[4854],M_list[4855],M_list[4856],M_list[4857],M_list[4858],M_list[4859],M_list[4860],M_list[4861],M_list[4862],M_list[4863],M_list[4864],M_list[4865],M_list[4866],M_list[4867],M_list[4868],M_list[4869],M_list[4870],M_list[4871],M_list[4872],M_list[4873],M_list[4874],M_list[4875],M_list[4876],M_list[4877],M_list[4878],M_list[4879],M_list[4880],M_list[4881],M_list[4882],M_list[4883],M_list[4884],M_list[4885],M_list[4886],M_list[4887],M_list[4888],M_list[4889],M_list[4890],M_list[4891],M_list[4892],M_list[4893],M_list[4894],M_list[4895],M_list[4896],M_list[4897],M_list[4898],M_list[4899],M_list[4900],M_list[4901],M_list[4902],M_list[4903],M_list[4904],M_list[4905],M_list[4906],M_list[4907],M_list[4908],M_list[4909],M_list[4910],M_list[4911],M_list[4912],M_list[4913],M_list[4914],M_list[4915],M_list[4916],M_list[4917],M_list[4918],M_list[4919],M_list[4920],M_list[4921],M_list[4922],M_list[4923],M_list[4924],M_list[4925],M_list[4926],M_list[4927],M_list[4928],M_list[4929],M_list[4930],M_list[4931],M_list[4932],M_list[4933],M_list[4934],M_list[4935],M_list[4936],M_list[4937],M_list[4938],M_list[4939],M_list[4940],M_list[4941],M_list[4942],M_list[4943],M_list[4944],M_list[4945],M_list[4946],M_list[4947],M_list[4948],M_list[4949],M_list[4950],M_list[4951],M_list[4952],M_list[4953],M_list[4954],M_list[4955],M_list[4956],M_list[4957],M_list[4958],M_list[4959],M_list[4960],M_list[4961],M_list[4962],M_list[4963],M_list[4964],M_list[4965],M_list[4966],M_list[4967],M_list[4968],M_list[4969],M_list[4970],M_list[4971],M_list[4972],M_list[4973],M_list[4974],M_list[4975],M_list[4976],M_list[4977],M_list[4978],M_list[4979],M_list[4980],M_list[4981],M_list[4982],M_list[4983],M_list[4984],M_list[4985],M_list[4986],M_list[4987],M_list[4988],M_list[4989],M_list[4990],M_list[4991],M_list[4992],M_list[4993],M_list[4994],M_list[4995],M_list[4996],M_list[4997],M_list[4998],M_list[4999],M_list[5000],M_list[5001],M_list[5002],M_list[5003],M_list[5004],M_list[5005],M_list[5006],M_list[5007],M_list[5008],M_list[5009],M_list[5010],M_list[5011],M_list[5012],M_list[5013],M_list[5014],M_list[5015],M_list[5016],M_list[5017],M_list[5018],M_list[5019],M_list[5020],M_list[5021],M_list[5022],M_list[5023],M_list[5024],M_list[5025],M_list[5026],M_list[5027],M_list[5028],M_list[5029],M_list[5030],M_list[5031],M_list[5032],M_list[5033],M_list[5034],M_list[5035],M_list[5036],M_list[5037],M_list[5038],M_list[5039],M_list[5040],M_list[5041],M_list[5042],M_list[5043],M_list[5044],M_list[5045],M_list[5046],M_list[5047],M_list[5048],M_list[5049],M_list[5050],M_list[5051],M_list[5052],M_list[5053],M_list[5054],M_list[5055],M_list[5056],M_list[5057],M_list[5058],M_list[5059],M_list[5060],M_list[5061],M_list[5062],M_list[5063],M_list[5064],M_list[5065],M_list[5066],M_list[5067],M_list[5068],M_list[5069],M_list[5070],M_list[5071],M_list[5072],M_list[5073],M_list[5074],M_list[5075],M_list[5076],M_list[5077],M_list[5078],M_list[5079],M_list[5080],M_list[5081],M_list[5082],M_list[5083],M_list[5084],M_list[5085],M_list[5086],M_list[5087],M_list[5088],M_list[5089],M_list[5090],M_list[5091],M_list[5092],M_list[5093],M_list[5094],M_list[5095],M_list[5096],M_list[5097],M_list[5098],M_list[5099],M_list[5100],M_list[5101],M_list[5102],M_list[5103],M_list[5104],M_list[5105],M_list[5106],M_list[5107],M_list[5108],M_list[5109],M_list[5110],M_list[5111],M_list[5112],M_list[5113],M_list[5114],M_list[5115],M_list[5116],M_list[5117],M_list[5118],M_list[5119],M_list[5120],M_list[5121],M_list[5122],M_list[5123],M_list[5124],M_list[5125],M_list[5126],M_list[5127],M_list[5128],M_list[5129],M_list[5130],M_list[5131],M_list[5132],M_list[5133],M_list[5134],M_list[5135],M_list[5136],M_list[5137],M_list[5138],M_list[5139],M_list[5140],M_list[5141],M_list[5142],M_list[5143],M_list[5144],M_list[5145],M_list[5146],M_list[5147],M_list[5148],M_list[5149],M_list[5150],M_list[5151],M_list[5152],M_list[5153],M_list[5154],M_list[5155],M_list[5156],M_list[5157],M_list[5158],M_list[5159],M_list[5160],M_list[5161],M_list[5162],M_list[5163],M_list[5164],M_list[5165],M_list[5166],M_list[5167],M_list[5168],M_list[5169],M_list[5170],M_list[5171],M_list[5172],M_list[5173],M_list[5174],M_list[5175],M_list[5176],M_list[5177],M_list[5178],M_list[5179],M_list[5180],M_list[5181],M_list[5182],M_list[5183],M_list[5184],M_list[5185],M_list[5186],M_list[5187],M_list[5188],M_list[5189],M_list[5190],M_list[5191],M_list[5192],M_list[5193],M_list[5194],M_list[5195],M_list[5196],M_list[5197],M_list[5198],M_list[5199],M_list[5200],M_list[5201],M_list[5202],M_list[5203],M_list[5204],M_list[5205],M_list[5206],M_list[5207],M_list[5208],M_list[5209],M_list[5210],M_list[5211],M_list[5212],M_list[5213],M_list[5214],M_list[5215],M_list[5216],M_list[5217],M_list[5218],M_list[5219],M_list[5220],M_list[5221],M_list[5222],M_list[5223],M_list[5224],M_list[5225],M_list[5226],M_list[5227],M_list[5228],M_list[5229],M_list[5230],M_list[5231],M_list[5232],M_list[5233],M_list[5234],M_list[5235],M_list[5236],M_list[5237],M_list[5238],M_list[5239],M_list[5240],M_list[5241],M_list[5242],M_list[5243],M_list[5244],M_list[5245],M_list[5246],M_list[5247],M_list[5248],M_list[5249],M_list[5250],M_list[5251],M_list[5252],M_list[5253],M_list[5254],M_list[5255],M_list[5256],M_list[5257],M_list[5258],M_list[5259],M_list[5260],M_list[5261],M_list[5262],M_list[5263],M_list[5264],M_list[5265],M_list[5266],M_list[5267],M_list[5268],M_list[5269],M_list[5270],M_list[5271],M_list[5272],M_list[5273],M_list[5274],M_list[5275],M_list[5276],M_list[5277],M_list[5278],M_list[5279],M_list[5280],M_list[5281],M_list[5282],M_list[5283],M_list[5284],M_list[5285],M_list[5286],M_list[5287],M_list[5288],M_list[5289],M_list[5290],M_list[5291],M_list[5292],M_list[5293],M_list[5294],M_list[5295],M_list[5296],M_list[5297],M_list[5298],M_list[5299],M_list[5300],M_list[5301],M_list[5302],M_list[5303],M_list[5304],M_list[5305],M_list[5306],M_list[5307],M_list[5308],M_list[5309],M_list[5310],M_list[5311],M_list[5312],M_list[5313],M_list[5314],M_list[5315],M_list[5316],M_list[5317],M_list[5318],M_list[5319],M_list[5320],M_list[5321],M_list[5322],M_list[5323],M_list[5324],M_list[5325],M_list[5326],M_list[5327],M_list[5328],M_list[5329],M_list[5330],M_list[5331],M_list[5332],M_list[5333],M_list[5334],M_list[5335],M_list[5336],M_list[5337],M_list[5338],M_list[5339],M_list[5340],M_list[5341],M_list[5342],M_list[5343],M_list[5344],M_list[5345],M_list[5346],M_list[5347],M_list[5348],M_list[5349],M_list[5350],M_list[5351],M_list[5352],M_list[5353],M_list[5354],M_list[5355],M_list[5356],M_list[5357],M_list[5358],M_list[5359],M_list[5360],M_list[5361],M_list[5362],M_list[5363],M_list[5364],M_list[5365],M_list[5366],M_list[5367],M_list[5368],M_list[5369],M_list[5370],M_list[5371],M_list[5372],M_list[5373],M_list[5374],M_list[5375],M_list[5376],M_list[5377],M_list[5378],M_list[5379],M_list[5380],M_list[5381],M_list[5382],M_list[5383],M_list[5384],M_list[5385],M_list[5386],M_list[5387],M_list[5388],M_list[5389],M_list[5390],M_list[5391],M_list[5392],M_list[5393],M_list[5394],M_list[5395],M_list[5396],M_list[5397],M_list[5398],M_list[5399],M_list[5400],M_list[5401],M_list[5402],M_list[5403],M_list[5404],M_list[5405],M_list[5406],M_list[5407],M_list[5408],M_list[5409],M_list[5410],M_list[5411],M_list[5412],M_list[5413],M_list[5414],M_list[5415],M_list[5416],M_list[5417],M_list[5418],M_list[5419],M_list[5420],M_list[5421],M_list[5422],M_list[5423],M_list[5424],M_list[5425],M_list[5426],M_list[5427],M_list[5428],M_list[5429],M_list[5430],M_list[5431],M_list[5432],M_list[5433],M_list[5434],M_list[5435],M_list[5436],M_list[5437],M_list[5438],M_list[5439],M_list[5440],M_list[5441],M_list[5442],M_list[5443],M_list[5444],M_list[5445],M_list[5446],M_list[5447],M_list[5448],M_list[5449],M_list[5450],M_list[5451],M_list[5452],M_list[5453],M_list[5454],M_list[5455],M_list[5456],M_list[5457],M_list[5458],M_list[5459],M_list[5460],M_list[5461],M_list[5462],M_list[5463],M_list[5464],M_list[5465],M_list[5466],M_list[5467],M_list[5468],M_list[5469],M_list[5470],M_list[5471],M_list[5472],M_list[5473],M_list[5474],M_list[5475],M_list[5476],M_list[5477],M_list[5478],M_list[5479],M_list[5480],M_list[5481],M_list[5482],M_list[5483],M_list[5484],M_list[5485],M_list[5486],M_list[5487],M_list[5488],M_list[5489],M_list[5490],M_list[5491],M_list[5492],M_list[5493],M_list[5494],M_list[5495],M_list[5496],M_list[5497],M_list[5498],M_list[5499],M_list[5500],M_list[5501],M_list[5502],M_list[5503],M_list[5504],M_list[5505],M_list[5506],M_list[5507],M_list[5508],M_list[5509],M_list[5510],M_list[5511],M_list[5512],M_list[5513],M_list[5514],M_list[5515],M_list[5516],M_list[5517],M_list[5518],M_list[5519],M_list[5520],M_list[5521],M_list[5522],M_list[5523],M_list[5524],M_list[5525],M_list[5526],M_list[5527],M_list[5528],M_list[5529],M_list[5530],M_list[5531],M_list[5532],M_list[5533],M_list[5534],M_list[5535],M_list[5536],M_list[5537],M_list[5538],M_list[5539],M_list[5540],M_list[5541],M_list[5542],M_list[5543],M_list[5544],M_list[5545],M_list[5546],M_list[5547],M_list[5548],M_list[5549],M_list[5550],M_list[5551],M_list[5552],M_list[5553],M_list[5554],M_list[5555],M_list[5556],M_list[5557],M_list[5558],M_list[5559],M_list[5560],M_list[5561],M_list[5562],M_list[5563],M_list[5564],M_list[5565],M_list[5566],M_list[5567],M_list[5568],M_list[5569],M_list[5570],M_list[5571],M_list[5572],M_list[5573],M_list[5574],M_list[5575],M_list[5576],M_list[5577],M_list[5578],M_list[5579],M_list[5580],M_list[5581],M_list[5582],M_list[5583],M_list[5584],M_list[5585],M_list[5586],M_list[5587],M_list[5588],M_list[5589],M_list[5590],M_list[5591],M_list[5592],M_list[5593],M_list[5594],M_list[5595],M_list[5596],M_list[5597],M_list[5598],M_list[5599],M_list[5600],M_list[5601],M_list[5602],M_list[5603],M_list[5604],M_list[5605],M_list[5606],M_list[5607],M_list[5608],M_list[5609],M_list[5610],M_list[5611],M_list[5612],M_list[5613],M_list[5614],M_list[5615],M_list[5616],M_list[5617],M_list[5618],M_list[5619],M_list[5620],M_list[5621],M_list[5622],M_list[5623],M_list[5624],M_list[5625],M_list[5626],M_list[5627],M_list[5628],M_list[5629],M_list[5630],M_list[5631],M_list[5632],M_list[5633],M_list[5634],M_list[5635],M_list[5636],M_list[5637],M_list[5638],M_list[5639],M_list[5640],M_list[5641],M_list[5642],M_list[5643],M_list[5644],M_list[5645],M_list[5646],M_list[5647],M_list[5648],M_list[5649],M_list[5650],M_list[5651],M_list[5652],M_list[5653],M_list[5654],M_list[5655],M_list[5656],M_list[5657],M_list[5658],M_list[5659],M_list[5660],M_list[5661],M_list[5662],M_list[5663],M_list[5664],M_list[5665],M_list[5666],M_list[5667],M_list[5668],M_list[5669],M_list[5670],M_list[5671],M_list[5672],M_list[5673],M_list[5674],M_list[5675],M_list[5676],M_list[5677],M_list[5678],M_list[5679],M_list[5680],M_list[5681],M_list[5682],M_list[5683],M_list[5684],M_list[5685],M_list[5686],M_list[5687],M_list[5688],M_list[5689],M_list[5690],M_list[5691],M_list[5692],M_list[5693],M_list[5694],M_list[5695],M_list[5696],M_list[5697],M_list[5698],M_list[5699],M_list[5700],M_list[5701],M_list[5702],M_list[5703],M_list[5704],M_list[5705],M_list[5706],M_list[5707],M_list[5708],M_list[5709],M_list[5710],M_list[5711],M_list[5712],M_list[5713],M_list[5714],M_list[5715],M_list[5716],M_list[5717],M_list[5718],M_list[5719],M_list[5720],M_list[5721],M_list[5722],M_list[5723],M_list[5724],M_list[5725],M_list[5726],M_list[5727],M_list[5728],M_list[5729],M_list[5730],M_list[5731],M_list[5732],M_list[5733],M_list[5734],M_list[5735],M_list[5736],M_list[5737],M_list[5738],M_list[5739],M_list[5740],M_list[5741],M_list[5742],M_list[5743],M_list[5744],M_list[5745],M_list[5746],M_list[5747],M_list[5748],M_list[5749],M_list[5750],M_list[5751],M_list[5752],M_list[5753],M_list[5754],M_list[5755],M_list[5756],M_list[5757],M_list[5758],M_list[5759],M_list[5760],M_list[5761],M_list[5762],M_list[5763],M_list[5764],M_list[5765],M_list[5766],M_list[5767],M_list[5768],M_list[5769],M_list[5770],M_list[5771],M_list[5772],M_list[5773],M_list[5774],M_list[5775],M_list[5776],M_list[5777],M_list[5778],M_list[5779],M_list[5780],M_list[5781],M_list[5782],M_list[5783],M_list[5784],M_list[5785],M_list[5786],M_list[5787],M_list[5788],M_list[5789],M_list[5790],M_list[5791],M_list[5792],M_list[5793],M_list[5794],M_list[5795],M_list[5796],M_list[5797],M_list[5798],M_list[5799],M_list[5800],M_list[5801],M_list[5802],M_list[5803],M_list[5804],M_list[5805],M_list[5806],M_list[5807],M_list[5808],M_list[5809],M_list[5810],M_list[5811],M_list[5812],M_list[5813],M_list[5814],M_list[5815],M_list[5816],M_list[5817],M_list[5818],M_list[5819],M_list[5820],M_list[5821],M_list[5822],M_list[5823],M_list[5824],M_list[5825],M_list[5826],M_list[5827],M_list[5828],M_list[5829],M_list[5830],M_list[5831],M_list[5832],M_list[5833],M_list[5834],M_list[5835],M_list[5836],M_list[5837],M_list[5838],M_list[5839],M_list[5840],M_list[5841],M_list[5842],M_list[5843],M_list[5844],M_list[5845],M_list[5846],M_list[5847],M_list[5848],M_list[5849],M_list[5850],M_list[5851],M_list[5852],M_list[5853],M_list[5854],M_list[5855],M_list[5856],M_list[5857],M_list[5858],M_list[5859],M_list[5860],M_list[5861],M_list[5862],M_list[5863],M_list[5864],M_list[5865],M_list[5866],M_list[5867],M_list[5868],M_list[5869],M_list[5870],M_list[5871],M_list[5872],M_list[5873],M_list[5874],M_list[5875],M_list[5876],M_list[5877],M_list[5878],M_list[5879],M_list[5880],M_list[5881],M_list[5882],M_list[5883],M_list[5884],M_list[5885],M_list[5886],M_list[5887],M_list[5888],M_list[5889],M_list[5890],M_list[5891],M_list[5892],M_list[5893],M_list[5894],M_list[5895],M_list[5896],M_list[5897],M_list[5898],M_list[5899],M_list[5900],M_list[5901],M_list[5902],M_list[5903],M_list[5904],M_list[5905],M_list[5906],M_list[5907],M_list[5908],M_list[5909],M_list[5910],M_list[5911],M_list[5912],M_list[5913],M_list[5914],M_list[5915],M_list[5916],M_list[5917],M_list[5918],M_list[5919],M_list[5920],M_list[5921],M_list[5922],M_list[5923],M_list[5924],M_list[5925],M_list[5926],M_list[5927],M_list[5928],M_list[5929],M_list[5930],M_list[5931],M_list[5932],M_list[5933],M_list[5934],M_list[5935],M_list[5936],M_list[5937],M_list[5938],M_list[5939],M_list[5940],M_list[5941],M_list[5942],M_list[5943],M_list[5944],M_list[5945],M_list[5946],M_list[5947],M_list[5948],M_list[5949],M_list[5950],M_list[5951],M_list[5952],M_list[5953],M_list[5954],M_list[5955],M_list[5956],M_list[5957],M_list[5958],M_list[5959],M_list[5960],M_list[5961],M_list[5962],M_list[5963],M_list[5964],M_list[5965],M_list[5966],M_list[5967],M_list[5968],M_list[5969],M_list[5970],M_list[5971],M_list[5972],M_list[5973],M_list[5974],M_list[5975],M_list[5976],M_list[5977],M_list[5978],M_list[5979],M_list[5980],M_list[5981],M_list[5982],M_list[5983],M_list[5984],M_list[5985],M_list[5986],M_list[5987],M_list[5988],M_list[5989],M_list[5990],M_list[5991],M_list[5992],M_list[5993],M_list[5994],M_list[5995],M_list[5996],M_list[5997],M_list[5998],M_list[5999],M_list[6000],M_list[6001],M_list[6002],M_list[6003],M_list[6004],M_list[6005],M_list[6006],M_list[6007],M_list[6008],M_list[6009],M_list[6010],M_list[6011],M_list[6012],M_list[6013],M_list[6014],M_list[6015],M_list[6016],M_list[6017],M_list[6018],M_list[6019],M_list[6020],M_list[6021],M_list[6022],M_list[6023],M_list[6024],M_list[6025],M_list[6026],M_list[6027],M_list[6028],M_list[6029],M_list[6030],M_list[6031],M_list[6032],M_list[6033],M_list[6034],M_list[6035],M_list[6036],M_list[6037],M_list[6038],M_list[6039],M_list[6040],M_list[6041],M_list[6042],M_list[6043],M_list[6044],M_list[6045],M_list[6046],M_list[6047],M_list[6048],M_list[6049],M_list[6050],M_list[6051],M_list[6052],M_list[6053],M_list[6054],M_list[6055],M_list[6056],M_list[6057],M_list[6058],M_list[6059],M_list[6060],M_list[6061],M_list[6062],M_list[6063],M_list[6064],M_list[6065],M_list[6066],M_list[6067],M_list[6068],M_list[6069],M_list[6070],M_list[6071],M_list[6072],M_list[6073],M_list[6074],M_list[6075],M_list[6076],M_list[6077],M_list[6078],M_list[6079],M_list[6080],M_list[6081],M_list[6082],M_list[6083],M_list[6084],M_list[6085],M_list[6086],M_list[6087],M_list[6088],M_list[6089],M_list[6090],M_list[6091],M_list[6092],M_list[6093],M_list[6094],M_list[6095],M_list[6096],M_list[6097],M_list[6098],M_list[6099],M_list[6100],M_list[6101],M_list[6102],M_list[6103],M_list[6104],M_list[6105],M_list[6106],M_list[6107],M_list[6108],M_list[6109],M_list[6110],M_list[6111],M_list[6112],M_list[6113],M_list[6114],M_list[6115],M_list[6116],M_list[6117],M_list[6118],M_list[6119],M_list[6120],M_list[6121],M_list[6122],M_list[6123],M_list[6124],M_list[6125],M_list[6126],M_list[6127],M_list[6128],M_list[6129],M_list[6130],M_list[6131],M_list[6132],M_list[6133],M_list[6134],M_list[6135],M_list[6136],M_list[6137],M_list[6138],M_list[6139],M_list[6140],M_list[6141],M_list[6142],M_list[6143],M_list[6144],M_list[6145],M_list[6146],M_list[6147],M_list[6148],M_list[6149],M_list[6150],M_list[6151],M_list[6152],M_list[6153],M_list[6154],M_list[6155],M_list[6156],M_list[6157],M_list[6158],M_list[6159],M_list[6160],M_list[6161],M_list[6162],M_list[6163],M_list[6164],M_list[6165],M_list[6166],M_list[6167],M_list[6168],M_list[6169],M_list[6170],M_list[6171],M_list[6172],M_list[6173],M_list[6174],M_list[6175],M_list[6176],M_list[6177],M_list[6178],M_list[6179],M_list[6180],M_list[6181],M_list[6182],M_list[6183],M_list[6184],M_list[6185],M_list[6186],M_list[6187],M_list[6188],M_list[6189],M_list[6190],M_list[6191],M_list[6192],M_list[6193],M_list[6194],M_list[6195],M_list[6196],M_list[6197],M_list[6198],M_list[6199],M_list[6200],M_list[6201],M_list[6202],M_list[6203],M_list[6204],M_list[6205],M_list[6206],M_list[6207],M_list[6208],M_list[6209],M_list[6210],M_list[6211],M_list[6212],M_list[6213],M_list[6214],M_list[6215],M_list[6216],M_list[6217],M_list[6218],M_list[6219],M_list[6220],M_list[6221],M_list[6222],M_list[6223],M_list[6224],M_list[6225],M_list[6226],M_list[6227],M_list[6228],M_list[6229],M_list[6230],M_list[6231],M_list[6232],M_list[6233],M_list[6234],M_list[6235],M_list[6236],M_list[6237],M_list[6238],M_list[6239],M_list[6240],M_list[6241],M_list[6242],M_list[6243],M_list[6244],M_list[6245],M_list[6246],M_list[6247],M_list[6248],M_list[6249],M_list[6250],M_list[6251],M_list[6252],M_list[6253],M_list[6254],M_list[6255],M_list[6256],M_list[6257],M_list[6258],M_list[6259],M_list[6260],M_list[6261],M_list[6262],M_list[6263],M_list[6264],M_list[6265],M_list[6266],M_list[6267],M_list[6268],M_list[6269],M_list[6270],M_list[6271],M_list[6272],M_list[6273],M_list[6274],M_list[6275],M_list[6276],M_list[6277],M_list[6278],M_list[6279],M_list[6280],M_list[6281],M_list[6282],M_list[6283],M_list[6284],M_list[6285],M_list[6286],M_list[6287],M_list[6288],M_list[6289],M_list[6290],M_list[6291],M_list[6292],M_list[6293],M_list[6294],M_list[6295],M_list[6296],M_list[6297],M_list[6298],M_list[6299],M_list[6300],M_list[6301],M_list[6302],M_list[6303],M_list[6304],M_list[6305],M_list[6306],M_list[6307],M_list[6308],M_list[6309],M_list[6310],M_list[6311],M_list[6312],M_list[6313],M_list[6314],M_list[6315],M_list[6316],M_list[6317],M_list[6318],M_list[6319],M_list[6320],M_list[6321],M_list[6322],M_list[6323],M_list[6324],M_list[6325],M_list[6326],M_list[6327],M_list[6328],M_list[6329],M_list[6330],M_list[6331],M_list[6332],M_list[6333],M_list[6334],M_list[6335],M_list[6336],M_list[6337],M_list[6338],M_list[6339],M_list[6340],M_list[6341],M_list[6342],M_list[6343],M_list[6344],M_list[6345],M_list[6346],M_list[6347],M_list[6348],M_list[6349],M_list[6350],M_list[6351],M_list[6352],M_list[6353],M_list[6354],M_list[6355],M_list[6356],M_list[6357],M_list[6358],M_list[6359],M_list[6360],M_list[6361],M_list[6362],M_list[6363],M_list[6364],M_list[6365],M_list[6366],M_list[6367],M_list[6368],M_list[6369],M_list[6370],M_list[6371],M_list[6372],M_list[6373],M_list[6374],M_list[6375],M_list[6376],M_list[6377],M_list[6378],M_list[6379],M_list[6380],M_list[6381],M_list[6382],M_list[6383],M_list[6384],M_list[6385],M_list[6386],M_list[6387],M_list[6388],M_list[6389],M_list[6390],M_list[6391],M_list[6392],M_list[6393],M_list[6394],M_list[6395],M_list[6396],M_list[6397],M_list[6398],M_list[6399]};

//pk 15
reg [7:0]pk_list[15:0];
wire [127:0]pk={pk_list[0],pk_list[1],pk_list[2],pk_list[3],pk_list[4],pk_list[5],pk_list[6],pk_list[7],pk_list[8],pk_list[9],pk_list[10],pk_list[11],pk_list[12],pk_list[13],pk_list[14],pk_list[15]};

reg [7:0]sk_list[15:0];
wire [127:0]sk={sk_list[0],sk_list[1],sk_list[2],sk_list[3],sk_list[4],sk_list[5],sk_list[6],sk_list[7],sk_list[8],sk_list[9],sk_list[10],sk_list[11],sk_list[12],sk_list[13],sk_list[14],sk_list[15]};


/*
module r_ram_for_verify
(
	input wire clk,
	input wire reset,
    input r_ram_for_verify_start,
	input [7:0] data, 


	output[14:0] address,
	output reg  r_ram_for_sign_end
);

//ht 31
wire [7:0]ht_list[31:0]

//salt 31
wire [7:0]salt_list[31:0]

//iSeedInfo 63
wire [7:0]iSeedInfo_list[63:0]

//cvInfo 127
wire [7:0]cvInfo_list[127:0]

//
//seedInfo 959
wire [7:0]seedInfo_list[959:0]

//masked_key 63
wire [7:0]masked_key_list[63:0]

//msgs 255
wire [7:0]msgs_list[255:0]

//C 127
wire [7:0]C_list[127:0]

//seed_lambda 255
wire [7:0]seed_lambda_list[255:0]

//aux_triangle 511
wire [7:0]aux_triangle_list[511:0]

// M 6399
wire [7:0]M_list[6399:0];

//pk 15
wire [7:0]pk_list[15:0]
*/

reg [14:0] counter1;  
reg [14:0] counter2;
reg counter3;
reg [5:0] state;

assign address=counter1;

reg signature_start;

wire signature_stop;

always @(posedge clk or negedge reset) begin
    if(~reset) begin
        r_ram_for_sign_end<=0;
        counter1<=0;
        counter2<=0;
        counter3<=0;
        state<=0;
        signature_start<=0;
    end
    else begin
        if(~r_ram_for_sign_start) begin
            r_ram_for_sign_end<=0;
            counter1<=0;
            counter2<=0;
            state<=0;
        end
        if(state==0&& r_ram_for_sign_start&&r_ram_for_sign_end==0) begin
            state<=1;
        end
        else if(state==1) begin
            if(~counter3) begin             
                counter1<=counter1+1;
                counter3<=~counter3;
            end
            else begin 
                counter3<=~counter3;
                if (counter2==6399) begin
                    counter2<=0;
                    state<=2;
                end
                else begin
                    counter2<=counter2+1;
                end
                M_list[counter2]<=data;
            end
        end
        else if(state==2) begin
            if(~counter3) begin             
                counter1<=counter1+1;
                counter3<=~counter3;
            end
            else begin 
                counter3<=~counter3;
                if (counter2==15) begin
                    counter2<=0;
                    state<=3;
                end
                else begin
                    counter2<=counter2+1;
                end
                pk_list[counter2]<=data;
            end
        end
        else if(state==3) begin
            if(~counter3) begin             
                counter1<=counter1+1;
                counter3<=~counter3;
            end
            else begin 
                counter3<=~counter3;
                if (counter2==15) begin
                    counter2<=0;
                    state<=4;
                end
                else begin
                    counter2<=counter2+1;
                end
                sk_list[counter2]<=data;
            end
        end
        else if(state==4) begin
            
            if(signature_stop==1) begin
                signature_start<=0;
                  state<=5;
            end
            else begin
                signature_start<=1;
            end
            
            //state<=5;
        end
        else if(state==5) begin
            counter1<=0;
            state<=0;
            r_ram_for_sign_end<=1;
        end
    end
end
/*
//ht 31
//salt 31
//iSeedInfo 63
//cvInfo 127
//seedInfo 959
//masked_key 63
//msgs 255
//C 127
//seed_lambda 255
//aux_triangle 511
//seed_triangle 15
// M 6399
//pk 15
*/
//assign sigma_out=M[19583:0];

sign_on_sm4_res1 sign(
    clk,
    reset,
    signature_start,
    M,
    sk,
    pk,
    signature_stop,
    sigma_out
);


endmodule 