`timescale 1ns / 1ps
/*
module testbench;
localparam
    CLK_FREQ    = 50_000_000,
    BAUD_RATE   = 115200,
    WORD_LENGTH = 8,
    STOP_BITS   = 2,
    PARITY      = "NONE";
reg clk, rst_n;
reg rx;
wire tx;

 top aa
(
				clk		,
				rst_n	,
				rx	,
				tx	
);


integer bitTime, idx, idxWord, idxBit;
reg [7:0] word [0:2];
reg [7:0]word2;
initial begin
    word2=2;
    clk = 0; rst_n = 0; rx = 1'b1; #10000; rst_n = 1; #10000;
    bitTime = 8680;  // ���ݲ���������λʱ������
    word[0] = 8'hfa; word[1] = 8'hff; word[2] = 8'ha5;
    for (idx=0; idx<10; idx=idx+1) begin  // �������
        for (idxWord=0; idxWord<1000000000; idxWord=idxWord+1) begin  // �����ֽ�
            rx = 1'b0; #bitTime; //start
            word2=0;
            for (idxBit=0; idxBit<8; idxBit=idxBit+1) begin  // ����λ
                rx = word2[idxBit];
                #bitTime;
            end
            rx = 1'b1; #bitTime; //stop
        end
        #1000000;
    end
end
always begin
    #10 clk = ~clk;
end
endmodule
*/

module tb();
    reg clk;
    reg reset;
    //input root_seed,
    //input salt
    reg sign_start;

    wire tapes;
     
     wire [255:0]H;
     wire [255:0]Cv;
     wire sign_end;
     wire verify_successful;
initial
begin
clk = 1'b0; 
reset = 1'b0; 

#100 reset = 1'b1; 
sign_start = 1'b1;

//data_i =1088'h0;
//#1000 wait(!sha3_busy) 
//h1InSeedSet[0:1087] =1088'h61616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161616161;
//h1InSeedSet[1088:1088*2-1]=0;
//h1InSeedSet[1088+1024]=1;
//h1InSeedSet[1088+59]=1;
//h1InSeedSet[1088+60]=1;
//h1InSeedSet[1088+61]=1;
//h1InSeedSet[1088+62]=1;
//h1InSeedSet[1088+63]=1;
wait(sign_end) sign_start =0;
wait(sign_end) sign_start =0;

end

wire verify_successful;

wire [255:0]Ht_i=256'h946544711A46346C513505B8DD4761F40B8B94A7577ED761376BD7A70F41190A;
wire [255:0]salt_i=256'h7D820E09EED566C7CC56D44802C4302E5C45D5B2B64B77391B0D21E1A60A4AD2;
wire [128*4-1:0]seed_star_i=512'h7953B1F113B617D6D9EBC3EB798344475D7BC112DD76530B7F29FBF5C843579FDEFE556178DC9418CA29AF4E3324D2519F822D3DB20CD54AD6EF3AE68C21FB00;
wire [256*4-1:0]Cv_i=1024'hCBDDE466EDF01BF5C1B8CB6260E707C14D166E54D9A973F0EA3C04FB97B7E42ACBDDE466EDF01BF5C1B8CB6260E707C14D166E54D9A973F0EA3C04FB97B7E42ACBDDE466EDF01BF5C1B8CB6260E707C14D166E54D9A973F0EA3C04FB97B7E42ACBDDE466EDF01BF5C1B8CB6260E707C14D166E54D9A973F0EA3C04FB97B7E42A;
wire [127:0] seed_triangle_i=128'h67B6E01D53F1CCCCD137EFFE087024E4;
wire [128*15*4-1:0]seedInfo=7680'hFA32714CF4EC5EFE934ABBFE482EC64839C2A3AC953701A596FEE0C8A3F78A520A9C8657D523ADEB87EA52566DB4842E2F1AFA2C90DD314B45CF363B77BA516456DC5A90C9084311FF03CDC15BBCECA29FC77B58D8C578D09229DD07B7A86FEF0E76F32D54863F5818623AB3EB8E76B03FC62BE4E0E2F928D34E7A3CD8007AD2A9D2FA7A3C876CBB15CB8F4F1C4ED997B1BF6569AF4B4FE76BA7FD56889C52BA4A23CCF9439F6F55FA0888B99F66D426D6776BEF267B3EDB1B9A55AA10947E5A47BE650C28D2686C9CC05F81DB3748D0DBAF8AADF19985661475F32F61B1BFC5EFA9DD5F2E17A3139F8EB1DF6E3B6F50DC5771EB6A85F7ED2ADAAC966FF9F57A56499336BA79C45B74DDAC18BE5975AC50ED708EC80032B7DF3274E7C7A404FB169466D70E520FCDCD77E8030B0201AF7D4B8781932FC1116C441949D0782FD698A06FD86E86352CCB36697B1FBCABF18089B9A2BE761A192D696A8A5330ABFB89BCFD29A986F862D20F54EA6F949B3C3CB0089DFCEA8DE30823760C0E71819D47E34262BC1CE9A3A9147E56CA1DF1953EB9A74A041DF7F9490FB3AD1EFD9AA704E9788654957C59EDCFB9432E79D4F47EDE9597351E5763F1650D7D5046CD18CEBE808C9B8BA8364B17724819166F93D71A2B01BF6C7E10791603F0D1AB8AF8FEC361E41ECDE2CA18A3FC201508B0B8DC5BF186A1E9F095C0E818356D067E1DEC83954A899E588264C7E2AA4DDBA21F7E58303452A89DDC8277453BD1AF707301A00CB30F0753AAFCC7FF25481162ECF6BE2C0F06C808B535038E04C472F8EF050974770B1D2A73FB339D5E7445638E34AB2ECCBD798C0F80FF632689BAB2F8A64BED3961649295E647690FF0D153BA4903594590D75590B5F5333B4D1926F01E343C305EAD425EFCC746B49BE47310C625E40644278CD1CB77EAA70DE8944EACA32C901EDAF2CBB781D5BC02DE8DB0E716C7E0EB85FDC5EDDCAB0E63103CFEDE2FE8D3A31C3815C8EB26043EFE39ECFF19F3875CAB28F01E78CE86050071EE8F15A8135115FC30E7EE978F13C0F406558EAAE4E4BE1C17664F82EA848ED8694B2CFF6BEBF8DF873DD362E44599B43BD82884C69684F4D8989C776C550A17F1182A4A4770DAE6BE231DA3BB6438679596C0B2AB3EA7B7218A95D4A669CDA36A7D46AF1FCA63AA48847CE24AF2B221ECA086DECD03B21EBB14B7AF54553950C8E73A252E2E84F598EFEC24CE1357FCC89ED239059D4CE2CFA10E50D637F585529BB90AD234607CC87E1F052F5A7D8B5724CF41C44EF58F83BADF9B0011B98A1B3B847A13C61F89CA18D6CB0FD6752F974B574BADEC8598275A9CC35C36F9D00C;
wire [128*4-1:0]masked_key=512'h7F1F3D434E86E8395CF2DFF02DE1EBC77F1F3D434E86E8395CF2DFF02DE1EBC77F1F3D434E86E8395CF2DFF02DE1EBC77F1F3D434E86E8395CF2DFF02DE1EBC7;
wire [512*4-1:0]msgs=2048'h8A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A79138A8A7913;
wire [256*4-1:0]C=1024'h1C68CA82A54DEADCA9F39CF2802ABB9C58610A83024B183B2EF14FE2F45C4B4EA1A3E383E765E92F9312A185DDACB45B4DC30C5F97DB29505151B8A127C2D0B501AFA737C35476483938A8F6872E7503B61DA1B5AFE61FA8B867B6DF2FEB9D3633C7057F762B3E3F6B53B6DD83E100618818871EE9D79AA0BBA23D0B74BBD3B3;
wire [512*4-1:0]seed_lambda=2048'h7DDBC6B11216C0C51DBC5359D227D5F6D44CE65D3BC3B55769C87BA6B3A0A23231347911A079EDB5D6DC85966EB38476CDC5B503D16AC0D6AC8A3093FA9617C656346959CF02D64226EB3B2EDC29BEC222E312E7ECE4374BC4FAB5760A698EEC770423C155791ED8F769AC62C8C55FC83FFA184CF18F4DB6A97B8BAA30EE20C63645B6C2DE769B73D8F334AF1AD68EB6BEEB0E9E4CC78CE9BFFB100B94733A106B4F9B4A97B6D96B5BDE06546F8CC3E63BF6CF71A69A73330CED73D4FCE46D64D17895472E2160E9B9BCE5C11F02FFB1D644337A77FAF63207B26A93388F4B343488BAE8FDA715CC8A43210940D92349C2D8B6ACC5FFE577D755E466E0BF543E;
wire [1024*4-1:0]aux_triangle=4096'h1C56458E1F8A4D17D3C9EBBE233C2802BA05A869975B3D14762475E76F9E2567D04BE8855519C8B50CEA63A8CE5418CEBC9A32C1C047C6FA7D15B08B0F9217C447ED96CF66C1EEC97D1C736B87E8A1F069F5BA9A63397E56AE134C061F012FBC32521B1EADA9ECE6CF144D786384361E222132657C3A430658CA02470DAE7C59EFA22A0443056918EE50B4489D7A45706DACC26EE2D360E18F229788C9332CF896A880BD57F04E8AE79E53CBCB1C723EB91C5EAEF04CAE56AAD818DF5869699492DDC8FE655D3EBE856F3155B61FDFBA9C81E105A2BAAC9F6CF8BC337111A77392445F9173EF6B3616605C25551687334D4C4A03DEEE786D021E65379AE001E16BC6375EC366F651156757EBCEFB55B052627917218668E5EF11F10B2FFF3BF094ECA15C717DE2DF28E62D38A5E723D9320BA1FDACFF417F09C0178D1A5AAE1852941C43261A20B8FC1C7C82CC91B65D56C63950AD75015FE8CE8FC893F0637F0302C5349764BF66B0F3073217B46811E033325B6FD828B045FC296706FA6F5ADA32647E07688808D8BE67677136738E7F595EAB22BD7B39C327DC5E5AF09D0BC934CC7E37BCF3487E85749985FFDEB91CD0D2C9C145D160790A982947507E075CA5E8A965B777829E34E4D173AF6BE70305184BE2330E0E350B20DADCB6F9AFEA2EDF8D79B47F20561A220E7E1A90D39AE5D1E1E70630758AB1EB183A1BA4CF;
 
    wire [51199:0]M=51200'h44463150407ceaee63ba0bfe5ad10d8f92705267f37682183cc8b29187fc7c4bdef3b892a413de80f8d726f59f112183d729ab4064e752b7c0b9c6053553b3e64f9f75f09f37a8720d77af0a312aaf1b4bc8f4c56aa772e3c7955ab6a7b179671e35160f5cd86e241563b965087fe4fbfe74a19509cb195d1cb9909a69b34b1897e9c71fdfd0f9f1322baa5ce997077d8ef7a40e4319f8974151b161f8f9163ffa795cbff955c29c2207e06389b0f582c17c79cce59df955d26d1597aac6d1c560839d57e99540c07a0002cd3319ef020b75d59952ed5aefce15cc617bfd3d9c3b2c0daff63ccea79b3667ee896eb1797054844d9a4378dfa1e50aa219ecb5532f5498d6252923f8f294b06eb223139039d62061d6d7796fea3940f43bce51fb898a42183793785b4bf22e7f4480ddd29483b598b71293effe01bd96bdfbe53d157c00a16f91c904d43bc7351eafc4e6790f0bf092e1ebd1034d87f04ff2782a6655be23bc3872f34e7384cd852de073819c4f13f240496bbe5e16b11e7c71e7d6608ed2d46eb9bbbeb64af2aba564b7cecedd8be5540f50dd0893c0a2c2775c15ed8ca705eeb6a1d0076d465a6a417e535ac2a76201945de652384def865247b45af6a2ac679b4b96adf140ae74376c7ee4f363a7fd2935af3c9d739725bc6728025b40778b076ab0b16a88b917fe14983f85fee06ebeee1dd7b6e1c00350ff16e1d7a014c3082b910f077a3982777a387d6c1206efa8c99f09d6d0706bff1399a9074a8cf1821e1bf1f20939dd65546cbc795d160ca9b2ddb70ca80c7792ea1cf7b9818f8abc8d7a3f09117e3bea233e47633d54c9fe0324e5b60b4fc0c82d61add9b3dab34e8bf36bd330047b77d79d83901c35cbd618ecd6f977ea3a30d2da56481d3a318b5ad70688d266559eed29ad36b38343ae97b99de0bb7d135f56ee67200999ad629c8f8d8caf2a41f944315645035ac599a75c06a996f2755b506eed32c856fbac883f048108c91f793b254ee42a9f63e675e02e8e5505b90179556bcd7ded1d8e792edb36293c3a106fbd33745b32ec95b8dc274e9a6c7a26540e5c2a145fcd8a5a9c8c77407ad4721bb7374f2dee807b629ff03cb450888ce7fd7c5b649e81d628a8936063cde5e665ae75035cd425ce317f1af6f722d183c62551ed7bd2eb2885da2d74b87912591273366a5167c21aff3ba34d8dac0948d2899e72fe62adebdc0745dd76a5e5a8e5047ada7edfcbedd9c3b5798555f7ccbab2f989fb382a6266f2687f7e3b98067cb01875ea218ca085deb9e2970ffbd1a471967bfd17e1e5e10a53fb0c4541108bc36c38de4f33d45f6f84d6774eb1b3bd81fa2f47b8ea81da9203d40e688f5a3d84303f37a230449ccaf4580fbed8a319d855ca4ed3009d4db01ced392d21fa84c5283633aeabd345cf94bea066fa1b794ed4bd15d522ee67f7f8292dbb245a9f0c981a386d742737af4e413b133351f253de9135a0800ff2361822d773c46f5eb4150132f4244718d8729877aa6048f72cdfb5bb6908a33d04044d02c09b37a72ca4e8317ee9b96a4a53b2c52b140f6db18c45c045f2932119313ac306d7acf814f7331dcbc51177a6a94e4cd12fab9fb38789b8711fb3b13ad460639ee668130b0dfc06291f0571750d8da7a0282ce38fc12f0175dd26c899898b0e4f4b1e458ef92848d2b06eea1a23dd1841deee9b3d4062ca97f5abd1460197e7ee712af04c5005df34a0f9d374023f5cfe469629aa0648fb90e7383ff3bcce7febd07d8ef0efa837ff99606ad9eba8540c1ef35b3912bcdf59a7d09a57806110dc868431000bdb6e0007298f3e838d3c1912a643585a846c27940bbcf867ed95de7f9ac939f3d410aca73f59dabb9aac0a6239538f33595a3879e5cced5d07f2b7c0944793240fd0e832e11420b7aec0b4180f7b6f8c1041c62e5261fad62162d7819537c75f788aebdef92bd55e9d9acbb4180b89706b2f4c199dd8ea975690aec9da370a19ee08027d18e46110b9bb86768e9ac66fbafcc1a4de2560d3f3628b2f39ce8028b98c1a13a684431dd906235b5b09b464e42d5e2930d4a3f509e71fae50990e5b1693cf75322f3f7ca11d3463eb040ecd2cb3a74d876902d755327e34fd7c7b2dc210b4f3c441974cc65482bc0ed7a7d5a62684595497d3a98c0d30664c5c7bc69194dc9db6789fa366b670bc725160946d5a2b7ea1a2b26dec420f2e33dac2115a37ce51aa3f7a903be4991bc03661247acbf76da9ce964ff75cbc32061f7a4ffead64c5352fd131e34d8b6460d050852e56a705fdd05c39c80a06068772c390b99ed0be6660ca61da0c7d22d42c430d047711b92903257d475f02f37811bf5c9caaa519a472047eb4a65dff5124d2f0bd7606099d1933798afde1dce311f638bf6c05152beec25b2bdb4ed918bb5587d97c5be9fffc55e6e85d8795c2cb03b74cd65fdf92409aa701dbebbfe4016ba05a7e25c74b183de36c82ad3aecbd4f46f7acddf9dd531f38cf9f5d950a901c1843c5f2fba5f638de8343bccee52ba3cba07f66df2f34422de9c0ec755614f283c51a51ab09e167da8aca2d52182636bbc350619b2ca4b325c9afbbddc676b08ae0e77332f56479088a99dfa829df5ab117764811950ffc19d03e5481757cef13ce93b55b49c5faed5c74562a4c2e64d47c1e5ddf97e6abed864232093357fa3dfe1e1b4e110bd414241d4a0ee63b969ed29f049e9855d24040a1467e59e328158ae17f822a2c1cc977d81288469d760a5c68612a3d7afffd3e2d85954ab501ed69ed380e74b46b4267d28c9c5c9034e61579cefd8110d4b788fb99ada93cef18c2c1c143a25bbdff3afec0edb0c30e42c6f5e985fe9a672a200ba5b04874c9c9798dfd45fc1911cda6ed0980faf394f559ab507454a5aebf64ece39b2f0f8f6806ddfeba1bd8dcd5c7fe8a7f058d01194818f461059b5d0ac00d8db679b21b4f11f7b0cdfb30728d3d3beb52803647f76401275fc1b37bbc9af17e7f38d407f6d5cef8676c7eb485bfd44cc07f157371d3d2894b362e959837019235ae73f5c14598a5fc639135ff3dc6920a04a6efb7ec89d3650f4e4547d3bd663e0ece84d351a32ebf00e60189831218c3b8a633db5068a561b934740651e1298eb1cf1c3fd0a2c642cfe92822629f615c8b38263a11f6b5cfd96b16a4e47bfa4d553add55cd8a11dcaca8c7fad49aebed8477c83df4fb272a4506a76660024ab86fe8212a739dc87f8d4f4c305a3ee6a153cfe30a12bdb1cbd707e7a5907aeb02569708a9349ee303b099e8be66ca6a7697b60d3c08293e956413841258de10d4b21ad52bb433655aa486ae9dd82991d0d12cefa95132d452472b375a8a16d17d87c142ba20c1b6b451bafeb48bca2c71f2256cfcf45cd028d3ce39b39749ef54255ed2ea5fba5a0e0ac397efc76c8b483695cce9c5415dde2e1873dd4fd7c4d93d50c4f0b1eb15cf12b8a9ba1f409b52e80f0cf10bdab8ee26042b62c0de72fb067735bac2104ab3e545328fda41d07767d2b0d828a90c2dad4bc12dc4300c801b850536edfae767e4c392696aa9bb8d281a15628926507828303a9e0037535c42c50e1b9d2ff136e9312e465c093af871abd7a47f458eafd1fc6b15feb5417955d536f57f74713c1f0a4779bbcab2981f472d36b9ffc394a5d687f615cdc6caa501f9c8fc8a49804dddc28f270c463447821d4ef940c3a15573af0d0942474d38cd82229697f1dcb3a07c4ca7b804fc91cfe2682ad52b2e22cd6f7bbabe469b2953296df8bb178a370bcc4347f6b38787dec13c4de162559f420553f62e42eab941cde6b9f4fc3be6719a90f91fe8042c3b108c9c6b4cf08a90497340c16dff3ac02d3889c3b987221c157aa71a285a946716ffcef0fac34b8dbb893e3250a18bc2a42fd3d71e76507d292716d184d3113146f0aceb7cf198a95ed07f698e556ef830054ca5773a29422840085d20cbba4e11a16edf874b135f80b227f13cddc5e910a201d0b81c36d68c9c441ffe34c243200b705090c69ef7eb4b832970f50d269341a10ccbccbf1b9fefb1ecfc426f6a179a2e6a3333e8e56ef23543f0dfdaa89ed8a92fec9e29da499b7f94a4f2e32c7a2fe396c3784e2313c76220eef9599f1d20fcfd21806ca6deca0ea0ae5efe786df408634458f183f5b8bec8d91487f798f2f7f607a03ca7cf0d11cdf14089c79e8ad82a7ab424fcf323b4429d52d3b04130bb657e667f2d72b9f0d558dd0e05b7d91cb013e8c8f119586887b3989da96089f967dd551590a80337f496922d0e2f25a2dc43eb69e951743f14feb241b6d02fada45b854248ce6b5469b7d344e7ef17e77ce3d1827a7c30498dca85e2540f948aa82e399c7c303e4637ec8ae4fbd624279b2c4e9eca6e137b1418192c42bb19d587e0a44b4fbf87e5a3a348f38f7e54169db07dfcada649ab2d98b0c8351a3f0f54c43c021b5c260dd99ef70e46036197fef3bac18af8430dba19407f17704aa2e8554e626982c0fd1efa32428aa7e0fabb263e750faa0d1f77686acc8b4e271a71f0010cdad9a60df718a7258d3d3c68d7aea2da8752e29b47abcb519ac21d4c9dbbe142ab5895b941b9a6082f452f48025c290153fc0cdcdf3e6dadcb7c6319dcf8f3ed59594af0e96d700972a2e60859b012c9c477872d614d0ccf45a61ee626a907f9bd8a53ca02da1eb9b84e5a198dc41125132f7c0b0ab389cbcec7f4ad0b9ac9a0f6a9350dcd44c84479fb23c4ee767813b6c794a63ce1f7bd2591552af09a6f12f477a99b5e2bf865375acb5f78f2dfeccc30ffa28f74997efae97f16f68f79a3ec72051a650b1928e5a8a6b910fbed10b181d02d20c7a81830d481cc723d5ae20658f358ad3a3c000b48d00d9e3ff9ec2dd0d9a2dac7b4502d735fdd00a600f4645ef43b49f1f51eb1c09be39051cf939a8bed55fc177e45ce744eb519b7dce5b46c9d22ca5828407de9dabae13b18871031cd0b12821a2e3d93ebb6a40823a87331fe5bc8d92dd04ac9020a0d2ccef39f86f347488c9bbc4be9a85723a8c26a992f72dd5611c6aaca6542b4a0129102b3c88c8e576bb37090b589d67a63ffed8bfcc03319b60098c7bfa3fb362b046f43718658bb2d410c9db6fbc3bfe27f1d04c781cd0d023404a3db58a6cce74457421d628541cc36edfd45dcd97aef15bf14a2117e54399500db5666b35d508391923f7c93cffbb8d320dd2a4f013bda7a571419e11f46e9fddeaaabce9351e72bc78a337255abeb083777411e877db66826b74ab7f28a9c26f8eab2386faa0239a3738f51fc9837179316ed038d0075934222bdce41611cfbcbb5632cf919d781c749395d6c1cbe2ce03d54ba82cb3156bb8de42b63450d7e79db69486e30855bc91b0546dee8536e697fb29f1cfa347e8c5d194befe09b29d35002aa21de23d755b481c43debdc47463400393ba3d5d9ab53dd698fe0f49eb224222dffd5b34cb10b5e5f181fce807e836b4dda5e04f1aae00d6695f93d1988b245b3bfa42e4c830ebb0c237ce60ec9e89dc82c05436a4ca858ab0d103b365d0d78b46d6438dff1d20ecdb1086a94aa62736e1966e9e1451888c7102a951f1834f7dd821b4eb8f88536676ca66707871520dfb4c7da390798a075152254c7da4a4eb297936acd4b18304069e54ed4b62f2a84e734c9a171f9a3ff44a54ab944884d6b89d2f50541a0a9565c00b7bd50cc553da8b693888a87fbac9edf03d4d6495c0b1258f2b870fc2794fabc82e1874d3f6f9bbf106bac304925d0ec768718f1eaef8e1f63fcc38d5a02306ed2c7562b6fc78265de731b06a8196626269fe135004e273a57ae68f249b8d731b0acbf0667b6f29c789f86af5b96577c92fe5d181d6ac8c8691226f79748d240b7555608044553da4c071b72fd3b77b50a7e6624955d366f84581ff97f02224d6d4ef949ce6d3454bf3921e6d89c820625e9ce3785af8edc89372001b79fa8412cd453981abaabc73c2ab67cdb2e73ce1da5dcf928f904f44921598d268a07463df5a0ad213727047fbee7eeea1223fe63e83f5558f31f01ef699abeb7f905d6f9bd142f7f9f5e320c16e0d36f1660eb62b42417a6f74d37d7aa9ea51ad1e340abdfd39d32d6e8d4f243a271859c46b8bf14768cb189bab3c54d63097f409244718d8c4ba9ae0c15609b788a1dc4130a427af3d0e17b515fe625186756aac4db06746b2e7cff0d3713fab71fa50321c3385c53817706385b516fff0d3584dbe8e602dba81d7c3296da1d65fa5bc06d8419dd7b26b8e49d713d1db8c5457e877175c5b7be0e7fbe7bfe42d11012ce5fdd4fc75783f3f05f488f19a324374f157a6fe8f6ca405bd2cfdf68c316e5bf9f710e555a135a25ffc075c62b9cd0426efd35101ca62a0e0f68651aa733bfca763c9c4b2867d459f2d163bef7f323217011d20975b4d1b302cbac753a0a5cbd49111f1414efb5b9609c979e14faaa74887ffbccff2ff145b68a44c7558e345a8778130a6c1f2de0c7fbbee9f795c87cfaf6db798df93cc2694609bedcd111bd68d44f4916dd7dd4e0c635906a6d2c3452f8ece14550d05406e0c8143b96095aa23a0d6b87dd89d10fddd545534dd91f324953b7300ac059bfb4955ddb34879a433c72c35ad91e62ebcb9ae378ed70b1723b34bcbcce7881831fe75e01bc5de08afa8981a419e549dffe62c01a1d0203b2f30a6b743c6d1a2e5fa95cc8dfc9d694eea89502a54f93247963c4f0078fb1aecef8632723693db51cdad514b97f157441ab383b54f044ab9f61d65c058d463f8808e4183d6cb83bda048ff18f693955055c0447cdbb773e6df1eb1249853b08d2fdce2824fb1c3eb2ab91c8e58c3444c2d23b4ddf875924dc1e371e6abd1866fa6b30aa252a7d9a5dcaa3ee73d3e695beb5a2439c9c35cfab2293fbe409538a6c6fe33bd7da3e76d56a6f052539251cae637ea4815ab46e643620477a9b6b9b00bcff74e7b07709931e67fb2251ab74c717f9d7391add70c6d023aa26905da84666baa4869a6f37da7d5d16fafbca952f9b2bd7ec5f74b1ae78080b5fea3f9036231d2704e4de9132df72376ef16819ce44e1a3a3ef982ce84367379d6d969df2000827405c072be3d1c4952e1a8edb0dff3553b1c9ddf77c6ecc7f27ed4973767b2ab982a15e933e384d95c35297f147b9f48480be2299c24669d66b4d52560b54295983712cdeff13db8c08677b6651a3298d586b442e637a3602b03454e95eaefa90c718d5be38642ea40fcf756646955cac7971b8344e396f12df2f527e08fd39e104fc13e14f90d2a1bbc580d68b4a15cda2955ef642e3b0e425ae8efd59a93e4324e629093ba5c779d69811e592c6482a1b393794771d1531624002c47004a50fe5fcfd7d646b1418930c3ebfed76646a2cfe70552ce4a3fd075c0b219ca752f5f371a10902c18e9396f530bd4d9416c56dc54ebef9d140f563eb0bd2fdf547e638fce723a502e637bbd1bd5bfc862fa07236c9ffc0afd2467432f8f5b1f1493c22c0ce7ba6d05d67116d639ddfdc3fab6137fba197a179e6b1dfb209169466c282e9f577d540b50426da8c07c1c37936dbf26678f0d0012ea6c90a3dfab2e60d1af237df9aaa4405622438602dbda8de380baeef2c7a48885b76e5b4e161facb47bbd756562e91776c86ad277b18d7eef0620a76fd111588bd18f2d36e689137ca673827d263327e628d55ba2e41f3a114165964b187a6f6cc049ad4165d493c77e9bb5198244d5e54fa872a617b88c784e14fbacc53b0098559e97f73687cd5c78f1f51de654dbfe9dd80aa6710ab705f66b9b186c525b315dbbaaead79a42ed3d66f491bd5e9e0abb62feb84e6728d5d026e42532ddbb375cac460e3fb8bdbb5497086d3665f2e08c43c9b0eb877e0ec386a905060520b079c3fa2b612eeec5325b9a01a47252936c9598ca3d649b9e1d429f54d0b857a28f539c4f523d436ca9c95e168e1d9fce7e3169f4ab80056466451ca78f2a409cd8d3153f6be8478db9947207685e1add3f45ee2bea131a25bc538d34d764d57ca63a29077ff13aa33d99d7832499c47a795722dc7fd25e4456614b55655cc61f80b7023b5ebf95f320e9e3740216a68faaaf4ca87bd937a6d7a710dc12fb2adc9e97276e239aec1902e877e5a131fa4dd38ed89e396000d81a45ee45012ca82227a2aba0afab3438371772cadd07438949e41197d433e1d53f48fe71235ce1fa9dec9ff50393eb8da93179550bf050c841830a6b89888fe526530861b56faaddb553db998cdd431b0d21c1ef5dc5010f1be07d2019ee359d149b996dfb4d4db7f00779358f0b0d232370947a6fe6562c0dcd5baebf47b0e49e51dae16536af7460b0610de2b502d7f05c1ede9e93d9955d7277143f3ee4a47c6d831ae3ffb0cd6f2065aac06e468f2fc44f34675abdb7fd9f14cfe32f2089400ef28b3e051e2e54c1a3c4bc70f865dd43dd026049e071663f05684ce0554e678e1f426710f3afbfcd486c97d38db48f29333631ee95c3af9fcefdc8fc86f900ab3dc2f0fa3bfc523104124d547a38f41eff44149efd850d14284c0456699ccbca5d07f4659b664954931023db1159aed96b741f1c86e9da20d192e7db7fdc2d8e037d372a0a3d97c9c9515a53b4919ed70b249fbd2e5d9f61c8e9048210c2f1e08dd3b4c10af95c6f78264d88a6c3c1b2580b2b1ab968d0ccfe685fe740df48e6bb67ce5a093a6475545a76fd7980519b7b7b3064d008dc8ca35fb52285b7872675c549411820065865f73a8e9846a5ac1c7e1b1352a8bc44537fef31d2dccc691452fe08cb93144f3226bfbc41e7af21d9128cd0ff30ec59418c02c734780761f1cfd911f47d6818fd8f21f722a4ec12f4cb424ef491b31e903f82f4856a948e16fb2d98a32eb1fc78e79ceb90f82520fcf5d948ab24f7b88cde50407ca938c6b4f79ab1d2bff964d460fe21e3ff58c42c72161e23536423373b4baaae0fc961af009766fa1086d4ba7e2fd410f;
    wire [127:0]pk=128'h0;


 verify_res1 vvv(
     clk,
     reset,
     8'h1,
    Ht_i,
    salt_i,
    seed_star_i,
    Cv_i,
    seed_triangle_i,
    //Z
   seedInfo,
    masked_key,
    msgs,
    C,
    seed_lambda,
   aux_triangle,

    M,
    pk,
     sign_start,
     H,
    verify_successful,
    sign_end
    );
    
always #5 clk = ~clk; //生成周期�????20ns，即频率�????50MHZ的时钟信号；


endmodule