module merkle_tree(
    input clk,
    input reset,
    //input c,
    //input salt
    input tree_start,
    output reg [511:0] commitment,
    output reg tree_set_end
    );
    wire[602*512-1:0] c=0;
    wire [0:255] salt=0;
    reg [1088-1:0] h3InCommitment [300:0];
    wire t=1;
    wire[15:0] j=1;
    wire [39:0]padding={8'h1f,24'h0,8'h80};
    wire [551:0]padding2={8'h1f,536'h0,8'h80};
    reg [300:0] Hstart;
    reg [300:0] restart;
    wire [511:0] hashValue[300:0];
    wire [300:0] en_end;
    wire [9:0] groupNum=1;
    reg[4:0] state; 
    reg[9:0] counter;
    wire [0:300] start_marsk[0:9];
    assign start_marsk[9] = 1;
    assign start_marsk[8] = 301'h3;
    assign start_marsk[7] = 301'h7;
    assign start_marsk[6] = 301'h1f;
    assign start_marsk[5] = 301'h3ff;
    assign start_marsk[4] = 301'h7ffff;
    assign start_marsk[3] = 301'h3fffffffff;
    assign start_marsk[2] = 301'hfffffffffffffffffff;
    assign start_marsk[1] = 301'h7fffffffffffffffffffffffffffffffffffff;
    assign start_marsk[0] = 301'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
    always @(posedge clk or negedge reset) begin
        if(~reset) begin
            counter <= 0;
            state<=0;
            tree_set_end<=0;
        end
        else begin
            if(state==0) begin
                if(tree_start) begin
                    tree_set_end<=0;
                    Hstart<=start_marsk[counter];
                    restart<=0;
                    state<=1;
                    if(counter==0)begin
                        h3InCommitment[0]={8'h03,c[308223:307712],c[307711:307200],j,padding};
                        h3InCommitment[1]={8'h03,c[307199:306688],c[306687:306176],j,padding};
                        h3InCommitment[2]={8'h03,c[306175:305664],c[305663:305152],j,padding};
                        h3InCommitment[3]={8'h03,c[305151:304640],c[304639:304128],j,padding};
                        h3InCommitment[4]={8'h03,c[304127:303616],c[303615:303104],j,padding};
                        h3InCommitment[5]={8'h03,c[303103:302592],c[302591:302080],j,padding};
                        h3InCommitment[6]={8'h03,c[302079:301568],c[301567:301056],j,padding};
                        h3InCommitment[7]={8'h03,c[301055:300544],c[300543:300032],j,padding};
                        h3InCommitment[8]={8'h03,c[300031:299520],c[299519:299008],j,padding};
                        h3InCommitment[9]={8'h03,c[299007:298496],c[298495:297984],j,padding};
                        h3InCommitment[10]={8'h03,c[297983:297472],c[297471:296960],j,padding};
                        h3InCommitment[11]={8'h03,c[296959:296448],c[296447:295936],j,padding};
                        h3InCommitment[12]={8'h03,c[295935:295424],c[295423:294912],j,padding};
                        h3InCommitment[13]={8'h03,c[294911:294400],c[294399:293888],j,padding};
                        h3InCommitment[14]={8'h03,c[293887:293376],c[293375:292864],j,padding};
                        h3InCommitment[15]={8'h03,c[292863:292352],c[292351:291840],j,padding};
                        h3InCommitment[16]={8'h03,c[291839:291328],c[291327:290816],j,padding};
                        h3InCommitment[17]={8'h03,c[290815:290304],c[290303:289792],j,padding};
                        h3InCommitment[18]={8'h03,c[289791:289280],c[289279:288768],j,padding};
                        h3InCommitment[19]={8'h03,c[288767:288256],c[288255:287744],j,padding};
                        h3InCommitment[20]={8'h03,c[287743:287232],c[287231:286720],j,padding};
                        h3InCommitment[21]={8'h03,c[286719:286208],c[286207:285696],j,padding};
                        h3InCommitment[22]={8'h03,c[285695:285184],c[285183:284672],j,padding};
                        h3InCommitment[23]={8'h03,c[284671:284160],c[284159:283648],j,padding};
                        h3InCommitment[24]={8'h03,c[283647:283136],c[283135:282624],j,padding};
                        h3InCommitment[25]={8'h03,c[282623:282112],c[282111:281600],j,padding};
                        h3InCommitment[26]={8'h03,c[281599:281088],c[281087:280576],j,padding};
                        h3InCommitment[27]={8'h03,c[280575:280064],c[280063:279552],j,padding};
                        h3InCommitment[28]={8'h03,c[279551:279040],c[279039:278528],j,padding};
                        h3InCommitment[29]={8'h03,c[278527:278016],c[278015:277504],j,padding};
                        h3InCommitment[30]={8'h03,c[277503:276992],c[276991:276480],j,padding};
                        h3InCommitment[31]={8'h03,c[276479:275968],c[275967:275456],j,padding};
                        h3InCommitment[32]={8'h03,c[275455:274944],c[274943:274432],j,padding};
                        h3InCommitment[33]={8'h03,c[274431:273920],c[273919:273408],j,padding};
                        h3InCommitment[34]={8'h03,c[273407:272896],c[272895:272384],j,padding};
                        h3InCommitment[35]={8'h03,c[272383:271872],c[271871:271360],j,padding};
                        h3InCommitment[36]={8'h03,c[271359:270848],c[270847:270336],j,padding};
                        h3InCommitment[37]={8'h03,c[270335:269824],c[269823:269312],j,padding};
                        h3InCommitment[38]={8'h03,c[269311:268800],c[268799:268288],j,padding};
                        h3InCommitment[39]={8'h03,c[268287:267776],c[267775:267264],j,padding};
                        h3InCommitment[40]={8'h03,c[267263:266752],c[266751:266240],j,padding};
                        h3InCommitment[41]={8'h03,c[266239:265728],c[265727:265216],j,padding};
                        h3InCommitment[42]={8'h03,c[265215:264704],c[264703:264192],j,padding};
                        h3InCommitment[43]={8'h03,c[264191:263680],c[263679:263168],j,padding};
                        h3InCommitment[44]={8'h03,c[263167:262656],c[262655:262144],j,padding};
                        h3InCommitment[45]={8'h03,c[262143:261632],c[261631:261120],j,padding};
                        h3InCommitment[46]={8'h03,c[261119:260608],c[260607:260096],j,padding};
                        h3InCommitment[47]={8'h03,c[260095:259584],c[259583:259072],j,padding};
                        h3InCommitment[48]={8'h03,c[259071:258560],c[258559:258048],j,padding};
                        h3InCommitment[49]={8'h03,c[258047:257536],c[257535:257024],j,padding};
                        h3InCommitment[50]={8'h03,c[257023:256512],c[256511:256000],j,padding};
                        h3InCommitment[51]={8'h03,c[255999:255488],c[255487:254976],j,padding};
                        h3InCommitment[52]={8'h03,c[254975:254464],c[254463:253952],j,padding};
                        h3InCommitment[53]={8'h03,c[253951:253440],c[253439:252928],j,padding};
                        h3InCommitment[54]={8'h03,c[252927:252416],c[252415:251904],j,padding};
                        h3InCommitment[55]={8'h03,c[251903:251392],c[251391:250880],j,padding};
                        h3InCommitment[56]={8'h03,c[250879:250368],c[250367:249856],j,padding};
                        h3InCommitment[57]={8'h03,c[249855:249344],c[249343:248832],j,padding};
                        h3InCommitment[58]={8'h03,c[248831:248320],c[248319:247808],j,padding};
                        h3InCommitment[59]={8'h03,c[247807:247296],c[247295:246784],j,padding};
                        h3InCommitment[60]={8'h03,c[246783:246272],c[246271:245760],j,padding};
                        h3InCommitment[61]={8'h03,c[245759:245248],c[245247:244736],j,padding};
                        h3InCommitment[62]={8'h03,c[244735:244224],c[244223:243712],j,padding};
                        h3InCommitment[63]={8'h03,c[243711:243200],c[243199:242688],j,padding};
                        h3InCommitment[64]={8'h03,c[242687:242176],c[242175:241664],j,padding};
                        h3InCommitment[65]={8'h03,c[241663:241152],c[241151:240640],j,padding};
                        h3InCommitment[66]={8'h03,c[240639:240128],c[240127:239616],j,padding};
                        h3InCommitment[67]={8'h03,c[239615:239104],c[239103:238592],j,padding};
                        h3InCommitment[68]={8'h03,c[238591:238080],c[238079:237568],j,padding};
                        h3InCommitment[69]={8'h03,c[237567:237056],c[237055:236544],j,padding};
                        h3InCommitment[70]={8'h03,c[236543:236032],c[236031:235520],j,padding};
                        h3InCommitment[71]={8'h03,c[235519:235008],c[235007:234496],j,padding};
                        h3InCommitment[72]={8'h03,c[234495:233984],c[233983:233472],j,padding};
                        h3InCommitment[73]={8'h03,c[233471:232960],c[232959:232448],j,padding};
                        h3InCommitment[74]={8'h03,c[232447:231936],c[231935:231424],j,padding};
                        h3InCommitment[75]={8'h03,c[231423:230912],c[230911:230400],j,padding};
                        h3InCommitment[76]={8'h03,c[230399:229888],c[229887:229376],j,padding};
                        h3InCommitment[77]={8'h03,c[229375:228864],c[228863:228352],j,padding};
                        h3InCommitment[78]={8'h03,c[228351:227840],c[227839:227328],j,padding};
                        h3InCommitment[79]={8'h03,c[227327:226816],c[226815:226304],j,padding};
                        h3InCommitment[80]={8'h03,c[226303:225792],c[225791:225280],j,padding};
                        h3InCommitment[81]={8'h03,c[225279:224768],c[224767:224256],j,padding};
                        h3InCommitment[82]={8'h03,c[224255:223744],c[223743:223232],j,padding};
                        h3InCommitment[83]={8'h03,c[223231:222720],c[222719:222208],j,padding};
                        h3InCommitment[84]={8'h03,c[222207:221696],c[221695:221184],j,padding};
                        h3InCommitment[85]={8'h03,c[221183:220672],c[220671:220160],j,padding};
                        h3InCommitment[86]={8'h03,c[220159:219648],c[219647:219136],j,padding};
                        h3InCommitment[87]={8'h03,c[219135:218624],c[218623:218112],j,padding};
                        h3InCommitment[88]={8'h03,c[218111:217600],c[217599:217088],j,padding};
                        h3InCommitment[89]={8'h03,c[217087:216576],c[216575:216064],j,padding};
                        h3InCommitment[90]={8'h03,c[216063:215552],c[215551:215040],j,padding};
                        h3InCommitment[91]={8'h03,c[215039:214528],c[214527:214016],j,padding};
                        h3InCommitment[92]={8'h03,c[214015:213504],c[213503:212992],j,padding};
                        h3InCommitment[93]={8'h03,c[212991:212480],c[212479:211968],j,padding};
                        h3InCommitment[94]={8'h03,c[211967:211456],c[211455:210944],j,padding};
                        h3InCommitment[95]={8'h03,c[210943:210432],c[210431:209920],j,padding};
                        h3InCommitment[96]={8'h03,c[209919:209408],c[209407:208896],j,padding};
                        h3InCommitment[97]={8'h03,c[208895:208384],c[208383:207872],j,padding};
                        h3InCommitment[98]={8'h03,c[207871:207360],c[207359:206848],j,padding};
                        h3InCommitment[99]={8'h03,c[206847:206336],c[206335:205824],j,padding};
                        h3InCommitment[100]={8'h03,c[205823:205312],c[205311:204800],j,padding};
                        h3InCommitment[101]={8'h03,c[204799:204288],c[204287:203776],j,padding};
                        h3InCommitment[102]={8'h03,c[203775:203264],c[203263:202752],j,padding};
                        h3InCommitment[103]={8'h03,c[202751:202240],c[202239:201728],j,padding};
                        h3InCommitment[104]={8'h03,c[201727:201216],c[201215:200704],j,padding};
                        h3InCommitment[105]={8'h03,c[200703:200192],c[200191:199680],j,padding};
                        h3InCommitment[106]={8'h03,c[199679:199168],c[199167:198656],j,padding};
                        h3InCommitment[107]={8'h03,c[198655:198144],c[198143:197632],j,padding};
                        h3InCommitment[108]={8'h03,c[197631:197120],c[197119:196608],j,padding};
                        h3InCommitment[109]={8'h03,c[196607:196096],c[196095:195584],j,padding};
                        h3InCommitment[110]={8'h03,c[195583:195072],c[195071:194560],j,padding};
                        h3InCommitment[111]={8'h03,c[194559:194048],c[194047:193536],j,padding};
                        h3InCommitment[112]={8'h03,c[193535:193024],c[193023:192512],j,padding};
                        h3InCommitment[113]={8'h03,c[192511:192000],c[191999:191488],j,padding};
                        h3InCommitment[114]={8'h03,c[191487:190976],c[190975:190464],j,padding};
                        h3InCommitment[115]={8'h03,c[190463:189952],c[189951:189440],j,padding};
                        h3InCommitment[116]={8'h03,c[189439:188928],c[188927:188416],j,padding};
                        h3InCommitment[117]={8'h03,c[188415:187904],c[187903:187392],j,padding};
                        h3InCommitment[118]={8'h03,c[187391:186880],c[186879:186368],j,padding};
                        h3InCommitment[119]={8'h03,c[186367:185856],c[185855:185344],j,padding};
                        h3InCommitment[120]={8'h03,c[185343:184832],c[184831:184320],j,padding};
                        h3InCommitment[121]={8'h03,c[184319:183808],c[183807:183296],j,padding};
                        h3InCommitment[122]={8'h03,c[183295:182784],c[182783:182272],j,padding};
                        h3InCommitment[123]={8'h03,c[182271:181760],c[181759:181248],j,padding};
                        h3InCommitment[124]={8'h03,c[181247:180736],c[180735:180224],j,padding};
                        h3InCommitment[125]={8'h03,c[180223:179712],c[179711:179200],j,padding};
                        h3InCommitment[126]={8'h03,c[179199:178688],c[178687:178176],j,padding};
                        h3InCommitment[127]={8'h03,c[178175:177664],c[177663:177152],j,padding};
                        h3InCommitment[128]={8'h03,c[177151:176640],c[176639:176128],j,padding};
                        h3InCommitment[129]={8'h03,c[176127:175616],c[175615:175104],j,padding};
                        h3InCommitment[130]={8'h03,c[175103:174592],c[174591:174080],j,padding};
                        h3InCommitment[131]={8'h03,c[174079:173568],c[173567:173056],j,padding};
                        h3InCommitment[132]={8'h03,c[173055:172544],c[172543:172032],j,padding};
                        h3InCommitment[133]={8'h03,c[172031:171520],c[171519:171008],j,padding};
                        h3InCommitment[134]={8'h03,c[171007:170496],c[170495:169984],j,padding};
                        h3InCommitment[135]={8'h03,c[169983:169472],c[169471:168960],j,padding};
                        h3InCommitment[136]={8'h03,c[168959:168448],c[168447:167936],j,padding};
                        h3InCommitment[137]={8'h03,c[167935:167424],c[167423:166912],j,padding};
                        h3InCommitment[138]={8'h03,c[166911:166400],c[166399:165888],j,padding};
                        h3InCommitment[139]={8'h03,c[165887:165376],c[165375:164864],j,padding};
                        h3InCommitment[140]={8'h03,c[164863:164352],c[164351:163840],j,padding};
                        h3InCommitment[141]={8'h03,c[163839:163328],c[163327:162816],j,padding};
                        h3InCommitment[142]={8'h03,c[162815:162304],c[162303:161792],j,padding};
                        h3InCommitment[143]={8'h03,c[161791:161280],c[161279:160768],j,padding};
                        h3InCommitment[144]={8'h03,c[160767:160256],c[160255:159744],j,padding};
                        h3InCommitment[145]={8'h03,c[159743:159232],c[159231:158720],j,padding};
                        h3InCommitment[146]={8'h03,c[158719:158208],c[158207:157696],j,padding};
                        h3InCommitment[147]={8'h03,c[157695:157184],c[157183:156672],j,padding};
                        h3InCommitment[148]={8'h03,c[156671:156160],c[156159:155648],j,padding};
                        h3InCommitment[149]={8'h03,c[155647:155136],c[155135:154624],j,padding};
                        h3InCommitment[150]={8'h03,c[154623:154112],c[154111:153600],j,padding};
                        h3InCommitment[151]={8'h03,c[153599:153088],c[153087:152576],j,padding};
                        h3InCommitment[152]={8'h03,c[152575:152064],c[152063:151552],j,padding};
                        h3InCommitment[153]={8'h03,c[151551:151040],c[151039:150528],j,padding};
                        h3InCommitment[154]={8'h03,c[150527:150016],c[150015:149504],j,padding};
                        h3InCommitment[155]={8'h03,c[149503:148992],c[148991:148480],j,padding};
                        h3InCommitment[156]={8'h03,c[148479:147968],c[147967:147456],j,padding};
                        h3InCommitment[157]={8'h03,c[147455:146944],c[146943:146432],j,padding};
                        h3InCommitment[158]={8'h03,c[146431:145920],c[145919:145408],j,padding};
                        h3InCommitment[159]={8'h03,c[145407:144896],c[144895:144384],j,padding};
                        h3InCommitment[160]={8'h03,c[144383:143872],c[143871:143360],j,padding};
                        h3InCommitment[161]={8'h03,c[143359:142848],c[142847:142336],j,padding};
                        h3InCommitment[162]={8'h03,c[142335:141824],c[141823:141312],j,padding};
                        h3InCommitment[163]={8'h03,c[141311:140800],c[140799:140288],j,padding};
                        h3InCommitment[164]={8'h03,c[140287:139776],c[139775:139264],j,padding};
                        h3InCommitment[165]={8'h03,c[139263:138752],c[138751:138240],j,padding};
                        h3InCommitment[166]={8'h03,c[138239:137728],c[137727:137216],j,padding};
                        h3InCommitment[167]={8'h03,c[137215:136704],c[136703:136192],j,padding};
                        h3InCommitment[168]={8'h03,c[136191:135680],c[135679:135168],j,padding};
                        h3InCommitment[169]={8'h03,c[135167:134656],c[134655:134144],j,padding};
                        h3InCommitment[170]={8'h03,c[134143:133632],c[133631:133120],j,padding};
                        h3InCommitment[171]={8'h03,c[133119:132608],c[132607:132096],j,padding};
                        h3InCommitment[172]={8'h03,c[132095:131584],c[131583:131072],j,padding};
                        h3InCommitment[173]={8'h03,c[131071:130560],c[130559:130048],j,padding};
                        h3InCommitment[174]={8'h03,c[130047:129536],c[129535:129024],j,padding};
                        h3InCommitment[175]={8'h03,c[129023:128512],c[128511:128000],j,padding};
                        h3InCommitment[176]={8'h03,c[127999:127488],c[127487:126976],j,padding};
                        h3InCommitment[177]={8'h03,c[126975:126464],c[126463:125952],j,padding};
                        h3InCommitment[178]={8'h03,c[125951:125440],c[125439:124928],j,padding};
                        h3InCommitment[179]={8'h03,c[124927:124416],c[124415:123904],j,padding};
                        h3InCommitment[180]={8'h03,c[123903:123392],c[123391:122880],j,padding};
                        h3InCommitment[181]={8'h03,c[122879:122368],c[122367:121856],j,padding};
                        h3InCommitment[182]={8'h03,c[121855:121344],c[121343:120832],j,padding};
                        h3InCommitment[183]={8'h03,c[120831:120320],c[120319:119808],j,padding};
                        h3InCommitment[184]={8'h03,c[119807:119296],c[119295:118784],j,padding};
                        h3InCommitment[185]={8'h03,c[118783:118272],c[118271:117760],j,padding};
                        h3InCommitment[186]={8'h03,c[117759:117248],c[117247:116736],j,padding};
                        h3InCommitment[187]={8'h03,c[116735:116224],c[116223:115712],j,padding};
                        h3InCommitment[188]={8'h03,c[115711:115200],c[115199:114688],j,padding};
                        h3InCommitment[189]={8'h03,c[114687:114176],c[114175:113664],j,padding};
                        h3InCommitment[190]={8'h03,c[113663:113152],c[113151:112640],j,padding};
                        h3InCommitment[191]={8'h03,c[112639:112128],c[112127:111616],j,padding};
                        h3InCommitment[192]={8'h03,c[111615:111104],c[111103:110592],j,padding};
                        h3InCommitment[193]={8'h03,c[110591:110080],c[110079:109568],j,padding};
                        h3InCommitment[194]={8'h03,c[109567:109056],c[109055:108544],j,padding};
                        h3InCommitment[195]={8'h03,c[108543:108032],c[108031:107520],j,padding};
                        h3InCommitment[196]={8'h03,c[107519:107008],c[107007:106496],j,padding};
                        h3InCommitment[197]={8'h03,c[106495:105984],c[105983:105472],j,padding};
                        h3InCommitment[198]={8'h03,c[105471:104960],c[104959:104448],j,padding};
                        h3InCommitment[199]={8'h03,c[104447:103936],c[103935:103424],j,padding};
                        h3InCommitment[200]={8'h03,c[103423:102912],c[102911:102400],j,padding};
                        h3InCommitment[201]={8'h03,c[102399:101888],c[101887:101376],j,padding};
                        h3InCommitment[202]={8'h03,c[101375:100864],c[100863:100352],j,padding};
                        h3InCommitment[203]={8'h03,c[100351:99840],c[99839:99328],j,padding};
                        h3InCommitment[204]={8'h03,c[99327:98816],c[98815:98304],j,padding};
                        h3InCommitment[205]={8'h03,c[98303:97792],c[97791:97280],j,padding};
                        h3InCommitment[206]={8'h03,c[97279:96768],c[96767:96256],j,padding};
                        h3InCommitment[207]={8'h03,c[96255:95744],c[95743:95232],j,padding};
                        h3InCommitment[208]={8'h03,c[95231:94720],c[94719:94208],j,padding};
                        h3InCommitment[209]={8'h03,c[94207:93696],c[93695:93184],j,padding};
                        h3InCommitment[210]={8'h03,c[93183:92672],c[92671:92160],j,padding};
                        h3InCommitment[211]={8'h03,c[92159:91648],c[91647:91136],j,padding};
                        h3InCommitment[212]={8'h03,c[91135:90624],c[90623:90112],j,padding};
                        h3InCommitment[213]={8'h03,c[90111:89600],c[89599:89088],j,padding};
                        h3InCommitment[214]={8'h03,c[89087:88576],c[88575:88064],j,padding};
                        h3InCommitment[215]={8'h03,c[88063:87552],c[87551:87040],j,padding};
                        h3InCommitment[216]={8'h03,c[87039:86528],c[86527:86016],j,padding};
                        h3InCommitment[217]={8'h03,c[86015:85504],c[85503:84992],j,padding};
                        h3InCommitment[218]={8'h03,c[84991:84480],c[84479:83968],j,padding};
                        h3InCommitment[219]={8'h03,c[83967:83456],c[83455:82944],j,padding};
                        h3InCommitment[220]={8'h03,c[82943:82432],c[82431:81920],j,padding};
                        h3InCommitment[221]={8'h03,c[81919:81408],c[81407:80896],j,padding};
                        h3InCommitment[222]={8'h03,c[80895:80384],c[80383:79872],j,padding};
                        h3InCommitment[223]={8'h03,c[79871:79360],c[79359:78848],j,padding};
                        h3InCommitment[224]={8'h03,c[78847:78336],c[78335:77824],j,padding};
                        h3InCommitment[225]={8'h03,c[77823:77312],c[77311:76800],j,padding};
                        h3InCommitment[226]={8'h03,c[76799:76288],c[76287:75776],j,padding};
                        h3InCommitment[227]={8'h03,c[75775:75264],c[75263:74752],j,padding};
                        h3InCommitment[228]={8'h03,c[74751:74240],c[74239:73728],j,padding};
                        h3InCommitment[229]={8'h03,c[73727:73216],c[73215:72704],j,padding};
                        h3InCommitment[230]={8'h03,c[72703:72192],c[72191:71680],j,padding};
                        h3InCommitment[231]={8'h03,c[71679:71168],c[71167:70656],j,padding};
                        h3InCommitment[232]={8'h03,c[70655:70144],c[70143:69632],j,padding};
                        h3InCommitment[233]={8'h03,c[69631:69120],c[69119:68608],j,padding};
                        h3InCommitment[234]={8'h03,c[68607:68096],c[68095:67584],j,padding};
                        h3InCommitment[235]={8'h03,c[67583:67072],c[67071:66560],j,padding};
                        h3InCommitment[236]={8'h03,c[66559:66048],c[66047:65536],j,padding};
                        h3InCommitment[237]={8'h03,c[65535:65024],c[65023:64512],j,padding};
                        h3InCommitment[238]={8'h03,c[64511:64000],c[63999:63488],j,padding};
                        h3InCommitment[239]={8'h03,c[63487:62976],c[62975:62464],j,padding};
                        h3InCommitment[240]={8'h03,c[62463:61952],c[61951:61440],j,padding};
                        h3InCommitment[241]={8'h03,c[61439:60928],c[60927:60416],j,padding};
                        h3InCommitment[242]={8'h03,c[60415:59904],c[59903:59392],j,padding};
                        h3InCommitment[243]={8'h03,c[59391:58880],c[58879:58368],j,padding};
                        h3InCommitment[244]={8'h03,c[58367:57856],c[57855:57344],j,padding};
                        h3InCommitment[245]={8'h03,c[57343:56832],c[56831:56320],j,padding};
                        h3InCommitment[246]={8'h03,c[56319:55808],c[55807:55296],j,padding};
                        h3InCommitment[247]={8'h03,c[55295:54784],c[54783:54272],j,padding};
                        h3InCommitment[248]={8'h03,c[54271:53760],c[53759:53248],j,padding};
                        h3InCommitment[249]={8'h03,c[53247:52736],c[52735:52224],j,padding};
                        h3InCommitment[250]={8'h03,c[52223:51712],c[51711:51200],j,padding};
                        h3InCommitment[251]={8'h03,c[51199:50688],c[50687:50176],j,padding};
                        h3InCommitment[252]={8'h03,c[50175:49664],c[49663:49152],j,padding};
                        h3InCommitment[253]={8'h03,c[49151:48640],c[48639:48128],j,padding};
                        h3InCommitment[254]={8'h03,c[48127:47616],c[47615:47104],j,padding};
                        h3InCommitment[255]={8'h03,c[47103:46592],c[46591:46080],j,padding};
                        h3InCommitment[256]={8'h03,c[46079:45568],c[45567:45056],j,padding};
                        h3InCommitment[257]={8'h03,c[45055:44544],c[44543:44032],j,padding};
                        h3InCommitment[258]={8'h03,c[44031:43520],c[43519:43008],j,padding};
                        h3InCommitment[259]={8'h03,c[43007:42496],c[42495:41984],j,padding};
                        h3InCommitment[260]={8'h03,c[41983:41472],c[41471:40960],j,padding};
                        h3InCommitment[261]={8'h03,c[40959:40448],c[40447:39936],j,padding};
                        h3InCommitment[262]={8'h03,c[39935:39424],c[39423:38912],j,padding};
                        h3InCommitment[263]={8'h03,c[38911:38400],c[38399:37888],j,padding};
                        h3InCommitment[264]={8'h03,c[37887:37376],c[37375:36864],j,padding};
                        h3InCommitment[265]={8'h03,c[36863:36352],c[36351:35840],j,padding};
                        h3InCommitment[266]={8'h03,c[35839:35328],c[35327:34816],j,padding};
                        h3InCommitment[267]={8'h03,c[34815:34304],c[34303:33792],j,padding};
                        h3InCommitment[268]={8'h03,c[33791:33280],c[33279:32768],j,padding};
                        h3InCommitment[269]={8'h03,c[32767:32256],c[32255:31744],j,padding};
                        h3InCommitment[270]={8'h03,c[31743:31232],c[31231:30720],j,padding};
                        h3InCommitment[271]={8'h03,c[30719:30208],c[30207:29696],j,padding};
                        h3InCommitment[272]={8'h03,c[29695:29184],c[29183:28672],j,padding};
                        h3InCommitment[273]={8'h03,c[28671:28160],c[28159:27648],j,padding};
                        h3InCommitment[274]={8'h03,c[27647:27136],c[27135:26624],j,padding};
                        h3InCommitment[275]={8'h03,c[26623:26112],c[26111:25600],j,padding};
                        h3InCommitment[276]={8'h03,c[25599:25088],c[25087:24576],j,padding};
                        h3InCommitment[277]={8'h03,c[24575:24064],c[24063:23552],j,padding};
                        h3InCommitment[278]={8'h03,c[23551:23040],c[23039:22528],j,padding};
                        h3InCommitment[279]={8'h03,c[22527:22016],c[22015:21504],j,padding};
                        h3InCommitment[280]={8'h03,c[21503:20992],c[20991:20480],j,padding};
                        h3InCommitment[281]={8'h03,c[20479:19968],c[19967:19456],j,padding};
                        h3InCommitment[282]={8'h03,c[19455:18944],c[18943:18432],j,padding};
                        h3InCommitment[283]={8'h03,c[18431:17920],c[17919:17408],j,padding};
                        h3InCommitment[284]={8'h03,c[17407:16896],c[16895:16384],j,padding};
                        h3InCommitment[285]={8'h03,c[16383:15872],c[15871:15360],j,padding};
                        h3InCommitment[286]={8'h03,c[15359:14848],c[14847:14336],j,padding};
                        h3InCommitment[287]={8'h03,c[14335:13824],c[13823:13312],j,padding};
                        h3InCommitment[288]={8'h03,c[13311:12800],c[12799:12288],j,padding};
                        h3InCommitment[289]={8'h03,c[12287:11776],c[11775:11264],j,padding};
                        h3InCommitment[290]={8'h03,c[11263:10752],c[10751:10240],j,padding};
                        h3InCommitment[291]={8'h03,c[10239:9728],c[9727:9216],j,padding};
                        h3InCommitment[292]={8'h03,c[9215:8704],c[8703:8192],j,padding};
                        h3InCommitment[293]={8'h03,c[8191:7680],c[7679:7168],j,padding};
                        h3InCommitment[294]={8'h03,c[7167:6656],c[6655:6144],j,padding};
                        h3InCommitment[295]={8'h03,c[6143:5632],c[5631:5120],j,padding};
                        h3InCommitment[296]={8'h03,c[5119:4608],c[4607:4096],j,padding};
                        h3InCommitment[297]={8'h03,c[4095:3584],c[3583:3072],j,padding};
                        h3InCommitment[298]={8'h03,c[3071:2560],c[2559:2048],j,padding};
                        h3InCommitment[299]={8'h03,c[2047:1536],c[1535:1024],j,padding};
                        h3InCommitment[300]={8'h03,c[1023:512],j,padding2};
                    end
                end
                
            end
            if(state==1) begin
                if(en_end==start_marsk[counter]) begin
                    counter<=counter+1;
                    restart<=Hstart;
                    if(en_end == start_marsk[9]) begin
                        state<=2;
                    end
                    else begin
                        state<=0;
                    end                        
                    h3InCommitment[0]<={8'h03,hashValue[0],hashValue[1],j,padding};
                    //h3InCommitment[1]<={8'h03,hashValue[2],hashValue[3],j,padding};
                    //h3InCommitment[2]<={8'h03,hashValue[4],hashValue[5],j,padding};
                    h3InCommitment[3]<={8'h03,hashValue[6],hashValue[7],j,padding};
                    h3InCommitment[4]<={8'h03,hashValue[8],hashValue[9],j,padding};
                    h3InCommitment[5]<={8'h03,hashValue[10],hashValue[11],j,padding};
                    h3InCommitment[6]<={8'h03,hashValue[12],hashValue[13],j,padding};
                    h3InCommitment[7]<={8'h03,hashValue[14],hashValue[15],j,padding};
                    h3InCommitment[8]<={8'h03,hashValue[16],hashValue[17],j,padding};
                    //h3InCommitment[9]<={8'h03,hashValue[18],hashValue[19],j,padding};
                    h3InCommitment[10]<={8'h03,hashValue[20],hashValue[21],j,padding};
                    h3InCommitment[11]<={8'h03,hashValue[22],hashValue[23],j,padding};
                    h3InCommitment[12]<={8'h03,hashValue[24],hashValue[25],j,padding};
                    h3InCommitment[13]<={8'h03,hashValue[26],hashValue[27],j,padding};
                    h3InCommitment[14]<={8'h03,hashValue[28],hashValue[29],j,padding};
                    h3InCommitment[15]<={8'h03,hashValue[30],hashValue[31],j,padding};
                    h3InCommitment[16]<={8'h03,hashValue[32],hashValue[33],j,padding};
                    h3InCommitment[17]<={8'h03,hashValue[34],hashValue[35],j,padding};
                    h3InCommitment[18]<={8'h03,hashValue[36],hashValue[37],j,padding};
                    h3InCommitment[19]<={8'h03,hashValue[38],hashValue[39],j,padding};
                    h3InCommitment[20]<={8'h03,hashValue[40],hashValue[41],j,padding};
                    h3InCommitment[21]<={8'h03,hashValue[42],hashValue[43],j,padding};
                    h3InCommitment[22]<={8'h03,hashValue[44],hashValue[45],j,padding};
                    h3InCommitment[23]<={8'h03,hashValue[46],hashValue[47],j,padding};
                    h3InCommitment[24]<={8'h03,hashValue[48],hashValue[49],j,padding};
                    h3InCommitment[25]<={8'h03,hashValue[50],hashValue[51],j,padding};
                    h3InCommitment[26]<={8'h03,hashValue[52],hashValue[53],j,padding};
                    h3InCommitment[27]<={8'h03,hashValue[54],hashValue[55],j,padding};
                    h3InCommitment[28]<={8'h03,hashValue[56],hashValue[57],j,padding};
                    h3InCommitment[29]<={8'h03,hashValue[58],hashValue[59],j,padding};
                    h3InCommitment[30]<={8'h03,hashValue[60],hashValue[61],j,padding};
                    h3InCommitment[31]<={8'h03,hashValue[62],hashValue[63],j,padding};
                    h3InCommitment[32]<={8'h03,hashValue[64],hashValue[65],j,padding};
                    h3InCommitment[33]<={8'h03,hashValue[66],hashValue[67],j,padding};
                    h3InCommitment[34]<={8'h03,hashValue[68],hashValue[69],j,padding};
                    h3InCommitment[35]<={8'h03,hashValue[70],hashValue[71],j,padding};
                    h3InCommitment[36]<={8'h03,hashValue[72],hashValue[73],j,padding};
                    h3InCommitment[37]<={8'h03,hashValue[74],hashValue[75],j,padding};
                    h3InCommitment[38]<={8'h03,hashValue[76],hashValue[77],j,padding};
                    h3InCommitment[39]<={8'h03,hashValue[78],hashValue[79],j,padding};
                    h3InCommitment[40]<={8'h03,hashValue[80],hashValue[81],j,padding};
                    h3InCommitment[41]<={8'h03,hashValue[82],hashValue[83],j,padding};
                    h3InCommitment[42]<={8'h03,hashValue[84],hashValue[85],j,padding};
                    h3InCommitment[43]<={8'h03,hashValue[86],hashValue[87],j,padding};
                    h3InCommitment[44]<={8'h03,hashValue[88],hashValue[89],j,padding};
                    h3InCommitment[45]<={8'h03,hashValue[90],hashValue[91],j,padding};
                    h3InCommitment[46]<={8'h03,hashValue[92],hashValue[93],j,padding};
                    h3InCommitment[47]<={8'h03,hashValue[94],hashValue[95],j,padding};
                    h3InCommitment[48]<={8'h03,hashValue[96],hashValue[97],j,padding};
                    h3InCommitment[49]<={8'h03,hashValue[98],hashValue[99],j,padding};
                    h3InCommitment[50]<={8'h03,hashValue[100],hashValue[101],j,padding};
                    h3InCommitment[51]<={8'h03,hashValue[102],hashValue[103],j,padding};
                    h3InCommitment[52]<={8'h03,hashValue[104],hashValue[105],j,padding};
                    h3InCommitment[53]<={8'h03,hashValue[106],hashValue[107],j,padding};
                    h3InCommitment[54]<={8'h03,hashValue[108],hashValue[109],j,padding};
                    h3InCommitment[55]<={8'h03,hashValue[110],hashValue[111],j,padding};
                    h3InCommitment[56]<={8'h03,hashValue[112],hashValue[113],j,padding};
                    h3InCommitment[57]<={8'h03,hashValue[114],hashValue[115],j,padding};
                    h3InCommitment[58]<={8'h03,hashValue[116],hashValue[117],j,padding};
                    h3InCommitment[59]<={8'h03,hashValue[118],hashValue[119],j,padding};
                    h3InCommitment[60]<={8'h03,hashValue[120],hashValue[121],j,padding};
                    h3InCommitment[61]<={8'h03,hashValue[122],hashValue[123],j,padding};
                    h3InCommitment[62]<={8'h03,hashValue[124],hashValue[125],j,padding};
                    h3InCommitment[63]<={8'h03,hashValue[126],hashValue[127],j,padding};
                    h3InCommitment[64]<={8'h03,hashValue[128],hashValue[129],j,padding};
                    h3InCommitment[65]<={8'h03,hashValue[130],hashValue[131],j,padding};
                    h3InCommitment[66]<={8'h03,hashValue[132],hashValue[133],j,padding};
                    h3InCommitment[67]<={8'h03,hashValue[134],hashValue[135],j,padding};
                    h3InCommitment[68]<={8'h03,hashValue[136],hashValue[137],j,padding};
                    h3InCommitment[69]<={8'h03,hashValue[138],hashValue[139],j,padding};
                    h3InCommitment[70]<={8'h03,hashValue[140],hashValue[141],j,padding};
                    h3InCommitment[71]<={8'h03,hashValue[142],hashValue[143],j,padding};
                    h3InCommitment[72]<={8'h03,hashValue[144],hashValue[145],j,padding};
                    h3InCommitment[73]<={8'h03,hashValue[146],hashValue[147],j,padding};
                    h3InCommitment[74]<={8'h03,hashValue[148],hashValue[149],j,padding};
                    //h3InCommitment[75]<={8'h03,hashValue[150],hashValue[151],j,padding};
                    h3InCommitment[76]<={8'h03,hashValue[152],hashValue[153],j,padding};
                    h3InCommitment[77]<={8'h03,hashValue[154],hashValue[155],j,padding};
                    h3InCommitment[78]<={8'h03,hashValue[156],hashValue[157],j,padding};
                    h3InCommitment[79]<={8'h03,hashValue[158],hashValue[159],j,padding};
                    h3InCommitment[80]<={8'h03,hashValue[160],hashValue[161],j,padding};
                    h3InCommitment[81]<={8'h03,hashValue[162],hashValue[163],j,padding};
                    h3InCommitment[82]<={8'h03,hashValue[164],hashValue[165],j,padding};
                    h3InCommitment[83]<={8'h03,hashValue[166],hashValue[167],j,padding};
                    h3InCommitment[84]<={8'h03,hashValue[168],hashValue[169],j,padding};
                    h3InCommitment[85]<={8'h03,hashValue[170],hashValue[171],j,padding};
                    h3InCommitment[86]<={8'h03,hashValue[172],hashValue[173],j,padding};
                    h3InCommitment[87]<={8'h03,hashValue[174],hashValue[175],j,padding};
                    h3InCommitment[88]<={8'h03,hashValue[176],hashValue[177],j,padding};
                    h3InCommitment[89]<={8'h03,hashValue[178],hashValue[179],j,padding};
                    h3InCommitment[90]<={8'h03,hashValue[180],hashValue[181],j,padding};
                    h3InCommitment[91]<={8'h03,hashValue[182],hashValue[183],j,padding};
                    h3InCommitment[92]<={8'h03,hashValue[184],hashValue[185],j,padding};
                    h3InCommitment[93]<={8'h03,hashValue[186],hashValue[187],j,padding};
                    h3InCommitment[94]<={8'h03,hashValue[188],hashValue[189],j,padding};
                    h3InCommitment[95]<={8'h03,hashValue[190],hashValue[191],j,padding};
                    h3InCommitment[96]<={8'h03,hashValue[192],hashValue[193],j,padding};
                    h3InCommitment[97]<={8'h03,hashValue[194],hashValue[195],j,padding};
                    h3InCommitment[98]<={8'h03,hashValue[196],hashValue[197],j,padding};
                    h3InCommitment[99]<={8'h03,hashValue[198],hashValue[199],j,padding};
                    h3InCommitment[100]<={8'h03,hashValue[200],hashValue[201],j,padding};
                    h3InCommitment[101]<={8'h03,hashValue[202],hashValue[203],j,padding};
                    h3InCommitment[102]<={8'h03,hashValue[204],hashValue[205],j,padding};
                    h3InCommitment[103]<={8'h03,hashValue[206],hashValue[207],j,padding};
                    h3InCommitment[104]<={8'h03,hashValue[208],hashValue[209],j,padding};
                    h3InCommitment[105]<={8'h03,hashValue[210],hashValue[211],j,padding};
                    h3InCommitment[106]<={8'h03,hashValue[212],hashValue[213],j,padding};
                    h3InCommitment[107]<={8'h03,hashValue[214],hashValue[215],j,padding};
                    h3InCommitment[108]<={8'h03,hashValue[216],hashValue[217],j,padding};
                    h3InCommitment[109]<={8'h03,hashValue[218],hashValue[219],j,padding};
                    h3InCommitment[110]<={8'h03,hashValue[220],hashValue[221],j,padding};
                    h3InCommitment[111]<={8'h03,hashValue[222],hashValue[223],j,padding};
                    h3InCommitment[112]<={8'h03,hashValue[224],hashValue[225],j,padding};
                    h3InCommitment[113]<={8'h03,hashValue[226],hashValue[227],j,padding};
                    h3InCommitment[114]<={8'h03,hashValue[228],hashValue[229],j,padding};
                    h3InCommitment[115]<={8'h03,hashValue[230],hashValue[231],j,padding};
                    h3InCommitment[116]<={8'h03,hashValue[232],hashValue[233],j,padding};
                    h3InCommitment[117]<={8'h03,hashValue[234],hashValue[235],j,padding};
                    h3InCommitment[118]<={8'h03,hashValue[236],hashValue[237],j,padding};
                    h3InCommitment[119]<={8'h03,hashValue[238],hashValue[239],j,padding};
                    h3InCommitment[120]<={8'h03,hashValue[240],hashValue[241],j,padding};
                    h3InCommitment[121]<={8'h03,hashValue[242],hashValue[243],j,padding};
                    h3InCommitment[122]<={8'h03,hashValue[244],hashValue[245],j,padding};
                    h3InCommitment[123]<={8'h03,hashValue[246],hashValue[247],j,padding};
                    h3InCommitment[124]<={8'h03,hashValue[248],hashValue[249],j,padding};
                    h3InCommitment[125]<={8'h03,hashValue[250],hashValue[251],j,padding};
                    h3InCommitment[126]<={8'h03,hashValue[252],hashValue[253],j,padding};
                    h3InCommitment[127]<={8'h03,hashValue[254],hashValue[255],j,padding};
                    h3InCommitment[128]<={8'h03,hashValue[256],hashValue[257],j,padding};
                    h3InCommitment[129]<={8'h03,hashValue[258],hashValue[259],j,padding};
                    h3InCommitment[130]<={8'h03,hashValue[260],hashValue[261],j,padding};
                    h3InCommitment[131]<={8'h03,hashValue[262],hashValue[263],j,padding};
                    h3InCommitment[132]<={8'h03,hashValue[264],hashValue[265],j,padding};
                    h3InCommitment[133]<={8'h03,hashValue[266],hashValue[267],j,padding};
                    h3InCommitment[134]<={8'h03,hashValue[268],hashValue[269],j,padding};
                    h3InCommitment[135]<={8'h03,hashValue[270],hashValue[271],j,padding};
                    h3InCommitment[136]<={8'h03,hashValue[272],hashValue[273],j,padding};
                    h3InCommitment[137]<={8'h03,hashValue[274],hashValue[275],j,padding};
                    h3InCommitment[138]<={8'h03,hashValue[276],hashValue[277],j,padding};
                    h3InCommitment[139]<={8'h03,hashValue[278],hashValue[279],j,padding};
                    h3InCommitment[140]<={8'h03,hashValue[280],hashValue[281],j,padding};
                    h3InCommitment[141]<={8'h03,hashValue[282],hashValue[283],j,padding};
                    h3InCommitment[142]<={8'h03,hashValue[284],hashValue[285],j,padding};
                    h3InCommitment[143]<={8'h03,hashValue[286],hashValue[287],j,padding};
                    h3InCommitment[144]<={8'h03,hashValue[288],hashValue[289],j,padding};
                    h3InCommitment[145]<={8'h03,hashValue[290],hashValue[291],j,padding};
                    h3InCommitment[146]<={8'h03,hashValue[292],hashValue[293],j,padding};
                    h3InCommitment[147]<={8'h03,hashValue[294],hashValue[295],j,padding};
                    h3InCommitment[148]<={8'h03,hashValue[296],hashValue[297],j,padding};
                    h3InCommitment[149]<={8'h03,hashValue[298],hashValue[299],j,padding};
                    h3InCommitment[150]<={8'h03,hashValue[300],j,padding2};
                    if(counter==2) begin
                        h3InCommitment[1]<={8'h03,hashValue[2],hashValue[3],j,padding};
                        h3InCommitment[2]<={8'h03,hashValue[4],hashValue[5],j,padding};
                        h3InCommitment[9]<={8'h03,hashValue[18],hashValue[19],j,padding};
                        h3InCommitment[75]<={8'h03,hashValue[150],j,padding2};
                    end
                    else if(counter==5) begin
                        h3InCommitment[1]<={8'h03,hashValue[2],hashValue[3],j,padding};
                        h3InCommitment[2]<={8'h03,hashValue[4],hashValue[5],j,padding};
                        h3InCommitment[9]<={8'h03,hashValue[18],j,padding2};
                    end
                    else if(counter==7) begin
                        h3InCommitment[1]<={8'h03,hashValue[2],hashValue[3],j,padding};
                        h3InCommitment[2]<={8'h03,hashValue[4],j,padding2};
                    end
                    else if(counter==8) begin
                        h3InCommitment[1]<={8'h03,hashValue[2],j,padding2};
                    end
                    else begin
                        h3InCommitment[1]<={8'h03,hashValue[2],hashValue[3],j,padding};
                        h3InCommitment[2]<={8'h03,hashValue[4],hashValue[5],j,padding};
                        h3InCommitment[9]<={8'h03,hashValue[18],hashValue[19],j,padding};
                        h3InCommitment[75]<={8'h03,hashValue[150],hashValue[151],j,padding};
                    end
                end
                                   
            end
            if(state==2) begin
                tree_set_end<=1;
                state <= 3;
            end
            if(state==3) begin
                tree_set_end <= 0;
                state<=0;
            end
        end

    end
    H h0(clk,reset,4'h1,2176'h0,h3InCommitment[0],Hstart[0],restart[0],groupNum,hashValue[0],en_end[0]);
    H h1(clk,reset,4'h1,2176'h0,h3InCommitment[1],Hstart[1],restart[1],groupNum,hashValue[1],en_end[1]);
    H h2(clk,reset,4'h1,2176'h0,h3InCommitment[2],Hstart[2],restart[2],groupNum,hashValue[2],en_end[2]);
    H h3(clk,reset,4'h1,2176'h0,h3InCommitment[3],Hstart[3],restart[3],groupNum,hashValue[3],en_end[3]);
    H h4(clk,reset,4'h1,2176'h0,h3InCommitment[4],Hstart[4],restart[4],groupNum,hashValue[4],en_end[4]);
    H h5(clk,reset,4'h1,2176'h0,h3InCommitment[5],Hstart[5],restart[5],groupNum,hashValue[5],en_end[5]);
    H h6(clk,reset,4'h1,2176'h0,h3InCommitment[6],Hstart[6],restart[6],groupNum,hashValue[6],en_end[6]);
    H h7(clk,reset,4'h1,2176'h0,h3InCommitment[7],Hstart[7],restart[7],groupNum,hashValue[7],en_end[7]);
    H h8(clk,reset,4'h1,2176'h0,h3InCommitment[8],Hstart[8],restart[8],groupNum,hashValue[8],en_end[8]);
    H h9(clk,reset,4'h1,2176'h0,h3InCommitment[9],Hstart[9],restart[9],groupNum,hashValue[9],en_end[9]);
    H h10(clk,reset,4'h1,2176'h0,h3InCommitment[10],Hstart[10],restart[10],groupNum,hashValue[10],en_end[10]);
    H h11(clk,reset,4'h1,2176'h0,h3InCommitment[11],Hstart[11],restart[11],groupNum,hashValue[11],en_end[11]);
    H h12(clk,reset,4'h1,2176'h0,h3InCommitment[12],Hstart[12],restart[12],groupNum,hashValue[12],en_end[12]);
    H h13(clk,reset,4'h1,2176'h0,h3InCommitment[13],Hstart[13],restart[13],groupNum,hashValue[13],en_end[13]);
    H h14(clk,reset,4'h1,2176'h0,h3InCommitment[14],Hstart[14],restart[14],groupNum,hashValue[14],en_end[14]);
    H h15(clk,reset,4'h1,2176'h0,h3InCommitment[15],Hstart[15],restart[15],groupNum,hashValue[15],en_end[15]);
    H h16(clk,reset,4'h1,2176'h0,h3InCommitment[16],Hstart[16],restart[16],groupNum,hashValue[16],en_end[16]);
    H h17(clk,reset,4'h1,2176'h0,h3InCommitment[17],Hstart[17],restart[17],groupNum,hashValue[17],en_end[17]);
    H h18(clk,reset,4'h1,2176'h0,h3InCommitment[18],Hstart[18],restart[18],groupNum,hashValue[18],en_end[18]);
    H h19(clk,reset,4'h1,2176'h0,h3InCommitment[19],Hstart[19],restart[19],groupNum,hashValue[19],en_end[19]);
    H h20(clk,reset,4'h1,2176'h0,h3InCommitment[20],Hstart[20],restart[20],groupNum,hashValue[20],en_end[20]);
    H h21(clk,reset,4'h1,2176'h0,h3InCommitment[21],Hstart[21],restart[21],groupNum,hashValue[21],en_end[21]);
    H h22(clk,reset,4'h1,2176'h0,h3InCommitment[22],Hstart[22],restart[22],groupNum,hashValue[22],en_end[22]);
    H h23(clk,reset,4'h1,2176'h0,h3InCommitment[23],Hstart[23],restart[23],groupNum,hashValue[23],en_end[23]);
    H h24(clk,reset,4'h1,2176'h0,h3InCommitment[24],Hstart[24],restart[24],groupNum,hashValue[24],en_end[24]);
    H h25(clk,reset,4'h1,2176'h0,h3InCommitment[25],Hstart[25],restart[25],groupNum,hashValue[25],en_end[25]);
    H h26(clk,reset,4'h1,2176'h0,h3InCommitment[26],Hstart[26],restart[26],groupNum,hashValue[26],en_end[26]);
    H h27(clk,reset,4'h1,2176'h0,h3InCommitment[27],Hstart[27],restart[27],groupNum,hashValue[27],en_end[27]);
    H h28(clk,reset,4'h1,2176'h0,h3InCommitment[28],Hstart[28],restart[28],groupNum,hashValue[28],en_end[28]);
    H h29(clk,reset,4'h1,2176'h0,h3InCommitment[29],Hstart[29],restart[29],groupNum,hashValue[29],en_end[29]);
    H h30(clk,reset,4'h1,2176'h0,h3InCommitment[30],Hstart[30],restart[30],groupNum,hashValue[30],en_end[30]);
    H h31(clk,reset,4'h1,2176'h0,h3InCommitment[31],Hstart[31],restart[31],groupNum,hashValue[31],en_end[31]);
    H h32(clk,reset,4'h1,2176'h0,h3InCommitment[32],Hstart[32],restart[32],groupNum,hashValue[32],en_end[32]);
    H h33(clk,reset,4'h1,2176'h0,h3InCommitment[33],Hstart[33],restart[33],groupNum,hashValue[33],en_end[33]);
    H h34(clk,reset,4'h1,2176'h0,h3InCommitment[34],Hstart[34],restart[34],groupNum,hashValue[34],en_end[34]);
    H h35(clk,reset,4'h1,2176'h0,h3InCommitment[35],Hstart[35],restart[35],groupNum,hashValue[35],en_end[35]);
    H h36(clk,reset,4'h1,2176'h0,h3InCommitment[36],Hstart[36],restart[36],groupNum,hashValue[36],en_end[36]);
    H h37(clk,reset,4'h1,2176'h0,h3InCommitment[37],Hstart[37],restart[37],groupNum,hashValue[37],en_end[37]);
    H h38(clk,reset,4'h1,2176'h0,h3InCommitment[38],Hstart[38],restart[38],groupNum,hashValue[38],en_end[38]);
    H h39(clk,reset,4'h1,2176'h0,h3InCommitment[39],Hstart[39],restart[39],groupNum,hashValue[39],en_end[39]);
    H h40(clk,reset,4'h1,2176'h0,h3InCommitment[40],Hstart[40],restart[40],groupNum,hashValue[40],en_end[40]);
    H h41(clk,reset,4'h1,2176'h0,h3InCommitment[41],Hstart[41],restart[41],groupNum,hashValue[41],en_end[41]);
    H h42(clk,reset,4'h1,2176'h0,h3InCommitment[42],Hstart[42],restart[42],groupNum,hashValue[42],en_end[42]);
    H h43(clk,reset,4'h1,2176'h0,h3InCommitment[43],Hstart[43],restart[43],groupNum,hashValue[43],en_end[43]);
    H h44(clk,reset,4'h1,2176'h0,h3InCommitment[44],Hstart[44],restart[44],groupNum,hashValue[44],en_end[44]);
    H h45(clk,reset,4'h1,2176'h0,h3InCommitment[45],Hstart[45],restart[45],groupNum,hashValue[45],en_end[45]);
    H h46(clk,reset,4'h1,2176'h0,h3InCommitment[46],Hstart[46],restart[46],groupNum,hashValue[46],en_end[46]);
    H h47(clk,reset,4'h1,2176'h0,h3InCommitment[47],Hstart[47],restart[47],groupNum,hashValue[47],en_end[47]);
    H h48(clk,reset,4'h1,2176'h0,h3InCommitment[48],Hstart[48],restart[48],groupNum,hashValue[48],en_end[48]);
    H h49(clk,reset,4'h1,2176'h0,h3InCommitment[49],Hstart[49],restart[49],groupNum,hashValue[49],en_end[49]);
    H h50(clk,reset,4'h1,2176'h0,h3InCommitment[50],Hstart[50],restart[50],groupNum,hashValue[50],en_end[50]);
    H h51(clk,reset,4'h1,2176'h0,h3InCommitment[51],Hstart[51],restart[51],groupNum,hashValue[51],en_end[51]);
    H h52(clk,reset,4'h1,2176'h0,h3InCommitment[52],Hstart[52],restart[52],groupNum,hashValue[52],en_end[52]);
    H h53(clk,reset,4'h1,2176'h0,h3InCommitment[53],Hstart[53],restart[53],groupNum,hashValue[53],en_end[53]);
    H h54(clk,reset,4'h1,2176'h0,h3InCommitment[54],Hstart[54],restart[54],groupNum,hashValue[54],en_end[54]);
    H h55(clk,reset,4'h1,2176'h0,h3InCommitment[55],Hstart[55],restart[55],groupNum,hashValue[55],en_end[55]);
    H h56(clk,reset,4'h1,2176'h0,h3InCommitment[56],Hstart[56],restart[56],groupNum,hashValue[56],en_end[56]);
    H h57(clk,reset,4'h1,2176'h0,h3InCommitment[57],Hstart[57],restart[57],groupNum,hashValue[57],en_end[57]);
    H h58(clk,reset,4'h1,2176'h0,h3InCommitment[58],Hstart[58],restart[58],groupNum,hashValue[58],en_end[58]);
    H h59(clk,reset,4'h1,2176'h0,h3InCommitment[59],Hstart[59],restart[59],groupNum,hashValue[59],en_end[59]);
    H h60(clk,reset,4'h1,2176'h0,h3InCommitment[60],Hstart[60],restart[60],groupNum,hashValue[60],en_end[60]);
    H h61(clk,reset,4'h1,2176'h0,h3InCommitment[61],Hstart[61],restart[61],groupNum,hashValue[61],en_end[61]);
    H h62(clk,reset,4'h1,2176'h0,h3InCommitment[62],Hstart[62],restart[62],groupNum,hashValue[62],en_end[62]);
    H h63(clk,reset,4'h1,2176'h0,h3InCommitment[63],Hstart[63],restart[63],groupNum,hashValue[63],en_end[63]);
    H h64(clk,reset,4'h1,2176'h0,h3InCommitment[64],Hstart[64],restart[64],groupNum,hashValue[64],en_end[64]);
    H h65(clk,reset,4'h1,2176'h0,h3InCommitment[65],Hstart[65],restart[65],groupNum,hashValue[65],en_end[65]);
    H h66(clk,reset,4'h1,2176'h0,h3InCommitment[66],Hstart[66],restart[66],groupNum,hashValue[66],en_end[66]);
    H h67(clk,reset,4'h1,2176'h0,h3InCommitment[67],Hstart[67],restart[67],groupNum,hashValue[67],en_end[67]);
    H h68(clk,reset,4'h1,2176'h0,h3InCommitment[68],Hstart[68],restart[68],groupNum,hashValue[68],en_end[68]);
    H h69(clk,reset,4'h1,2176'h0,h3InCommitment[69],Hstart[69],restart[69],groupNum,hashValue[69],en_end[69]);
    H h70(clk,reset,4'h1,2176'h0,h3InCommitment[70],Hstart[70],restart[70],groupNum,hashValue[70],en_end[70]);
    H h71(clk,reset,4'h1,2176'h0,h3InCommitment[71],Hstart[71],restart[71],groupNum,hashValue[71],en_end[71]);
    H h72(clk,reset,4'h1,2176'h0,h3InCommitment[72],Hstart[72],restart[72],groupNum,hashValue[72],en_end[72]);
    H h73(clk,reset,4'h1,2176'h0,h3InCommitment[73],Hstart[73],restart[73],groupNum,hashValue[73],en_end[73]);
    H h74(clk,reset,4'h1,2176'h0,h3InCommitment[74],Hstart[74],restart[74],groupNum,hashValue[74],en_end[74]);
    H h75(clk,reset,4'h1,2176'h0,h3InCommitment[75],Hstart[75],restart[75],groupNum,hashValue[75],en_end[75]);
    H h76(clk,reset,4'h1,2176'h0,h3InCommitment[76],Hstart[76],restart[76],groupNum,hashValue[76],en_end[76]);
    H h77(clk,reset,4'h1,2176'h0,h3InCommitment[77],Hstart[77],restart[77],groupNum,hashValue[77],en_end[77]);
    H h78(clk,reset,4'h1,2176'h0,h3InCommitment[78],Hstart[78],restart[78],groupNum,hashValue[78],en_end[78]);
    H h79(clk,reset,4'h1,2176'h0,h3InCommitment[79],Hstart[79],restart[79],groupNum,hashValue[79],en_end[79]);
    H h80(clk,reset,4'h1,2176'h0,h3InCommitment[80],Hstart[80],restart[80],groupNum,hashValue[80],en_end[80]);
    H h81(clk,reset,4'h1,2176'h0,h3InCommitment[81],Hstart[81],restart[81],groupNum,hashValue[81],en_end[81]);
    H h82(clk,reset,4'h1,2176'h0,h3InCommitment[82],Hstart[82],restart[82],groupNum,hashValue[82],en_end[82]);
    H h83(clk,reset,4'h1,2176'h0,h3InCommitment[83],Hstart[83],restart[83],groupNum,hashValue[83],en_end[83]);
    H h84(clk,reset,4'h1,2176'h0,h3InCommitment[84],Hstart[84],restart[84],groupNum,hashValue[84],en_end[84]);
    H h85(clk,reset,4'h1,2176'h0,h3InCommitment[85],Hstart[85],restart[85],groupNum,hashValue[85],en_end[85]);
    H h86(clk,reset,4'h1,2176'h0,h3InCommitment[86],Hstart[86],restart[86],groupNum,hashValue[86],en_end[86]);
    H h87(clk,reset,4'h1,2176'h0,h3InCommitment[87],Hstart[87],restart[87],groupNum,hashValue[87],en_end[87]);
    H h88(clk,reset,4'h1,2176'h0,h3InCommitment[88],Hstart[88],restart[88],groupNum,hashValue[88],en_end[88]);
    H h89(clk,reset,4'h1,2176'h0,h3InCommitment[89],Hstart[89],restart[89],groupNum,hashValue[89],en_end[89]);
    H h90(clk,reset,4'h1,2176'h0,h3InCommitment[90],Hstart[90],restart[90],groupNum,hashValue[90],en_end[90]);
    H h91(clk,reset,4'h1,2176'h0,h3InCommitment[91],Hstart[91],restart[91],groupNum,hashValue[91],en_end[91]);
    H h92(clk,reset,4'h1,2176'h0,h3InCommitment[92],Hstart[92],restart[92],groupNum,hashValue[92],en_end[92]);
    H h93(clk,reset,4'h1,2176'h0,h3InCommitment[93],Hstart[93],restart[93],groupNum,hashValue[93],en_end[93]);
    H h94(clk,reset,4'h1,2176'h0,h3InCommitment[94],Hstart[94],restart[94],groupNum,hashValue[94],en_end[94]);
    H h95(clk,reset,4'h1,2176'h0,h3InCommitment[95],Hstart[95],restart[95],groupNum,hashValue[95],en_end[95]);
    H h96(clk,reset,4'h1,2176'h0,h3InCommitment[96],Hstart[96],restart[96],groupNum,hashValue[96],en_end[96]);
    H h97(clk,reset,4'h1,2176'h0,h3InCommitment[97],Hstart[97],restart[97],groupNum,hashValue[97],en_end[97]);
    H h98(clk,reset,4'h1,2176'h0,h3InCommitment[98],Hstart[98],restart[98],groupNum,hashValue[98],en_end[98]);
    H h99(clk,reset,4'h1,2176'h0,h3InCommitment[99],Hstart[99],restart[99],groupNum,hashValue[99],en_end[99]);
    H h100(clk,reset,4'h1,2176'h0,h3InCommitment[100],Hstart[100],restart[100],groupNum,hashValue[100],en_end[100]);
    H h101(clk,reset,4'h1,2176'h0,h3InCommitment[101],Hstart[101],restart[101],groupNum,hashValue[101],en_end[101]);
    H h102(clk,reset,4'h1,2176'h0,h3InCommitment[102],Hstart[102],restart[102],groupNum,hashValue[102],en_end[102]);
    H h103(clk,reset,4'h1,2176'h0,h3InCommitment[103],Hstart[103],restart[103],groupNum,hashValue[103],en_end[103]);
    H h104(clk,reset,4'h1,2176'h0,h3InCommitment[104],Hstart[104],restart[104],groupNum,hashValue[104],en_end[104]);
    H h105(clk,reset,4'h1,2176'h0,h3InCommitment[105],Hstart[105],restart[105],groupNum,hashValue[105],en_end[105]);
    H h106(clk,reset,4'h1,2176'h0,h3InCommitment[106],Hstart[106],restart[106],groupNum,hashValue[106],en_end[106]);
    H h107(clk,reset,4'h1,2176'h0,h3InCommitment[107],Hstart[107],restart[107],groupNum,hashValue[107],en_end[107]);
    H h108(clk,reset,4'h1,2176'h0,h3InCommitment[108],Hstart[108],restart[108],groupNum,hashValue[108],en_end[108]);
    H h109(clk,reset,4'h1,2176'h0,h3InCommitment[109],Hstart[109],restart[109],groupNum,hashValue[109],en_end[109]);
    H h110(clk,reset,4'h1,2176'h0,h3InCommitment[110],Hstart[110],restart[110],groupNum,hashValue[110],en_end[110]);
    H h111(clk,reset,4'h1,2176'h0,h3InCommitment[111],Hstart[111],restart[111],groupNum,hashValue[111],en_end[111]);
    H h112(clk,reset,4'h1,2176'h0,h3InCommitment[112],Hstart[112],restart[112],groupNum,hashValue[112],en_end[112]);
    H h113(clk,reset,4'h1,2176'h0,h3InCommitment[113],Hstart[113],restart[113],groupNum,hashValue[113],en_end[113]);
    H h114(clk,reset,4'h1,2176'h0,h3InCommitment[114],Hstart[114],restart[114],groupNum,hashValue[114],en_end[114]);
    H h115(clk,reset,4'h1,2176'h0,h3InCommitment[115],Hstart[115],restart[115],groupNum,hashValue[115],en_end[115]);
    H h116(clk,reset,4'h1,2176'h0,h3InCommitment[116],Hstart[116],restart[116],groupNum,hashValue[116],en_end[116]);
    H h117(clk,reset,4'h1,2176'h0,h3InCommitment[117],Hstart[117],restart[117],groupNum,hashValue[117],en_end[117]);
    H h118(clk,reset,4'h1,2176'h0,h3InCommitment[118],Hstart[118],restart[118],groupNum,hashValue[118],en_end[118]);
    H h119(clk,reset,4'h1,2176'h0,h3InCommitment[119],Hstart[119],restart[119],groupNum,hashValue[119],en_end[119]);
    H h120(clk,reset,4'h1,2176'h0,h3InCommitment[120],Hstart[120],restart[120],groupNum,hashValue[120],en_end[120]);
    H h121(clk,reset,4'h1,2176'h0,h3InCommitment[121],Hstart[121],restart[121],groupNum,hashValue[121],en_end[121]);
    H h122(clk,reset,4'h1,2176'h0,h3InCommitment[122],Hstart[122],restart[122],groupNum,hashValue[122],en_end[122]);
    H h123(clk,reset,4'h1,2176'h0,h3InCommitment[123],Hstart[123],restart[123],groupNum,hashValue[123],en_end[123]);
    H h124(clk,reset,4'h1,2176'h0,h3InCommitment[124],Hstart[124],restart[124],groupNum,hashValue[124],en_end[124]);
    H h125(clk,reset,4'h1,2176'h0,h3InCommitment[125],Hstart[125],restart[125],groupNum,hashValue[125],en_end[125]);
    H h126(clk,reset,4'h1,2176'h0,h3InCommitment[126],Hstart[126],restart[126],groupNum,hashValue[126],en_end[126]);
    H h127(clk,reset,4'h1,2176'h0,h3InCommitment[127],Hstart[127],restart[127],groupNum,hashValue[127],en_end[127]);
    H h128(clk,reset,4'h1,2176'h0,h3InCommitment[128],Hstart[128],restart[128],groupNum,hashValue[128],en_end[128]);
    H h129(clk,reset,4'h1,2176'h0,h3InCommitment[129],Hstart[129],restart[129],groupNum,hashValue[129],en_end[129]);
    H h130(clk,reset,4'h1,2176'h0,h3InCommitment[130],Hstart[130],restart[130],groupNum,hashValue[130],en_end[130]);
    H h131(clk,reset,4'h1,2176'h0,h3InCommitment[131],Hstart[131],restart[131],groupNum,hashValue[131],en_end[131]);
    H h132(clk,reset,4'h1,2176'h0,h3InCommitment[132],Hstart[132],restart[132],groupNum,hashValue[132],en_end[132]);
    H h133(clk,reset,4'h1,2176'h0,h3InCommitment[133],Hstart[133],restart[133],groupNum,hashValue[133],en_end[133]);
    H h134(clk,reset,4'h1,2176'h0,h3InCommitment[134],Hstart[134],restart[134],groupNum,hashValue[134],en_end[134]);
    H h135(clk,reset,4'h1,2176'h0,h3InCommitment[135],Hstart[135],restart[135],groupNum,hashValue[135],en_end[135]);
    H h136(clk,reset,4'h1,2176'h0,h3InCommitment[136],Hstart[136],restart[136],groupNum,hashValue[136],en_end[136]);
    H h137(clk,reset,4'h1,2176'h0,h3InCommitment[137],Hstart[137],restart[137],groupNum,hashValue[137],en_end[137]);
    H h138(clk,reset,4'h1,2176'h0,h3InCommitment[138],Hstart[138],restart[138],groupNum,hashValue[138],en_end[138]);
    H h139(clk,reset,4'h1,2176'h0,h3InCommitment[139],Hstart[139],restart[139],groupNum,hashValue[139],en_end[139]);
    H h140(clk,reset,4'h1,2176'h0,h3InCommitment[140],Hstart[140],restart[140],groupNum,hashValue[140],en_end[140]);
    H h141(clk,reset,4'h1,2176'h0,h3InCommitment[141],Hstart[141],restart[141],groupNum,hashValue[141],en_end[141]);
    H h142(clk,reset,4'h1,2176'h0,h3InCommitment[142],Hstart[142],restart[142],groupNum,hashValue[142],en_end[142]);
    H h143(clk,reset,4'h1,2176'h0,h3InCommitment[143],Hstart[143],restart[143],groupNum,hashValue[143],en_end[143]);
    H h144(clk,reset,4'h1,2176'h0,h3InCommitment[144],Hstart[144],restart[144],groupNum,hashValue[144],en_end[144]);
    H h145(clk,reset,4'h1,2176'h0,h3InCommitment[145],Hstart[145],restart[145],groupNum,hashValue[145],en_end[145]);
    H h146(clk,reset,4'h1,2176'h0,h3InCommitment[146],Hstart[146],restart[146],groupNum,hashValue[146],en_end[146]);
    H h147(clk,reset,4'h1,2176'h0,h3InCommitment[147],Hstart[147],restart[147],groupNum,hashValue[147],en_end[147]);
    H h148(clk,reset,4'h1,2176'h0,h3InCommitment[148],Hstart[148],restart[148],groupNum,hashValue[148],en_end[148]);
    H h149(clk,reset,4'h1,2176'h0,h3InCommitment[149],Hstart[149],restart[149],groupNum,hashValue[149],en_end[149]);
    H h150(clk,reset,4'h1,2176'h0,h3InCommitment[150],Hstart[150],restart[150],groupNum,hashValue[150],en_end[150]);
    H h151(clk,reset,4'h1,2176'h0,h3InCommitment[151],Hstart[151],restart[151],groupNum,hashValue[151],en_end[151]);
    H h152(clk,reset,4'h1,2176'h0,h3InCommitment[152],Hstart[152],restart[152],groupNum,hashValue[152],en_end[152]);
    H h153(clk,reset,4'h1,2176'h0,h3InCommitment[153],Hstart[153],restart[153],groupNum,hashValue[153],en_end[153]);
    H h154(clk,reset,4'h1,2176'h0,h3InCommitment[154],Hstart[154],restart[154],groupNum,hashValue[154],en_end[154]);
    H h155(clk,reset,4'h1,2176'h0,h3InCommitment[155],Hstart[155],restart[155],groupNum,hashValue[155],en_end[155]);
    H h156(clk,reset,4'h1,2176'h0,h3InCommitment[156],Hstart[156],restart[156],groupNum,hashValue[156],en_end[156]);
    H h157(clk,reset,4'h1,2176'h0,h3InCommitment[157],Hstart[157],restart[157],groupNum,hashValue[157],en_end[157]);
    H h158(clk,reset,4'h1,2176'h0,h3InCommitment[158],Hstart[158],restart[158],groupNum,hashValue[158],en_end[158]);
    H h159(clk,reset,4'h1,2176'h0,h3InCommitment[159],Hstart[159],restart[159],groupNum,hashValue[159],en_end[159]);
    H h160(clk,reset,4'h1,2176'h0,h3InCommitment[160],Hstart[160],restart[160],groupNum,hashValue[160],en_end[160]);
    H h161(clk,reset,4'h1,2176'h0,h3InCommitment[161],Hstart[161],restart[161],groupNum,hashValue[161],en_end[161]);
    H h162(clk,reset,4'h1,2176'h0,h3InCommitment[162],Hstart[162],restart[162],groupNum,hashValue[162],en_end[162]);
    H h163(clk,reset,4'h1,2176'h0,h3InCommitment[163],Hstart[163],restart[163],groupNum,hashValue[163],en_end[163]);
    H h164(clk,reset,4'h1,2176'h0,h3InCommitment[164],Hstart[164],restart[164],groupNum,hashValue[164],en_end[164]);
    H h165(clk,reset,4'h1,2176'h0,h3InCommitment[165],Hstart[165],restart[165],groupNum,hashValue[165],en_end[165]);
    H h166(clk,reset,4'h1,2176'h0,h3InCommitment[166],Hstart[166],restart[166],groupNum,hashValue[166],en_end[166]);
    H h167(clk,reset,4'h1,2176'h0,h3InCommitment[167],Hstart[167],restart[167],groupNum,hashValue[167],en_end[167]);
    H h168(clk,reset,4'h1,2176'h0,h3InCommitment[168],Hstart[168],restart[168],groupNum,hashValue[168],en_end[168]);
    H h169(clk,reset,4'h1,2176'h0,h3InCommitment[169],Hstart[169],restart[169],groupNum,hashValue[169],en_end[169]);
    H h170(clk,reset,4'h1,2176'h0,h3InCommitment[170],Hstart[170],restart[170],groupNum,hashValue[170],en_end[170]);
    H h171(clk,reset,4'h1,2176'h0,h3InCommitment[171],Hstart[171],restart[171],groupNum,hashValue[171],en_end[171]);
    H h172(clk,reset,4'h1,2176'h0,h3InCommitment[172],Hstart[172],restart[172],groupNum,hashValue[172],en_end[172]);
    H h173(clk,reset,4'h1,2176'h0,h3InCommitment[173],Hstart[173],restart[173],groupNum,hashValue[173],en_end[173]);
    H h174(clk,reset,4'h1,2176'h0,h3InCommitment[174],Hstart[174],restart[174],groupNum,hashValue[174],en_end[174]);
    H h175(clk,reset,4'h1,2176'h0,h3InCommitment[175],Hstart[175],restart[175],groupNum,hashValue[175],en_end[175]);
    H h176(clk,reset,4'h1,2176'h0,h3InCommitment[176],Hstart[176],restart[176],groupNum,hashValue[176],en_end[176]);
    H h177(clk,reset,4'h1,2176'h0,h3InCommitment[177],Hstart[177],restart[177],groupNum,hashValue[177],en_end[177]);
    H h178(clk,reset,4'h1,2176'h0,h3InCommitment[178],Hstart[178],restart[178],groupNum,hashValue[178],en_end[178]);
    H h179(clk,reset,4'h1,2176'h0,h3InCommitment[179],Hstart[179],restart[179],groupNum,hashValue[179],en_end[179]);
    H h180(clk,reset,4'h1,2176'h0,h3InCommitment[180],Hstart[180],restart[180],groupNum,hashValue[180],en_end[180]);
    H h181(clk,reset,4'h1,2176'h0,h3InCommitment[181],Hstart[181],restart[181],groupNum,hashValue[181],en_end[181]);
    H h182(clk,reset,4'h1,2176'h0,h3InCommitment[182],Hstart[182],restart[182],groupNum,hashValue[182],en_end[182]);
    H h183(clk,reset,4'h1,2176'h0,h3InCommitment[183],Hstart[183],restart[183],groupNum,hashValue[183],en_end[183]);
    H h184(clk,reset,4'h1,2176'h0,h3InCommitment[184],Hstart[184],restart[184],groupNum,hashValue[184],en_end[184]);
    H h185(clk,reset,4'h1,2176'h0,h3InCommitment[185],Hstart[185],restart[185],groupNum,hashValue[185],en_end[185]);
    H h186(clk,reset,4'h1,2176'h0,h3InCommitment[186],Hstart[186],restart[186],groupNum,hashValue[186],en_end[186]);
    H h187(clk,reset,4'h1,2176'h0,h3InCommitment[187],Hstart[187],restart[187],groupNum,hashValue[187],en_end[187]);
    H h188(clk,reset,4'h1,2176'h0,h3InCommitment[188],Hstart[188],restart[188],groupNum,hashValue[188],en_end[188]);
    H h189(clk,reset,4'h1,2176'h0,h3InCommitment[189],Hstart[189],restart[189],groupNum,hashValue[189],en_end[189]);
    H h190(clk,reset,4'h1,2176'h0,h3InCommitment[190],Hstart[190],restart[190],groupNum,hashValue[190],en_end[190]);
    H h191(clk,reset,4'h1,2176'h0,h3InCommitment[191],Hstart[191],restart[191],groupNum,hashValue[191],en_end[191]);
    H h192(clk,reset,4'h1,2176'h0,h3InCommitment[192],Hstart[192],restart[192],groupNum,hashValue[192],en_end[192]);
    H h193(clk,reset,4'h1,2176'h0,h3InCommitment[193],Hstart[193],restart[193],groupNum,hashValue[193],en_end[193]);
    H h194(clk,reset,4'h1,2176'h0,h3InCommitment[194],Hstart[194],restart[194],groupNum,hashValue[194],en_end[194]);
    H h195(clk,reset,4'h1,2176'h0,h3InCommitment[195],Hstart[195],restart[195],groupNum,hashValue[195],en_end[195]);
    H h196(clk,reset,4'h1,2176'h0,h3InCommitment[196],Hstart[196],restart[196],groupNum,hashValue[196],en_end[196]);
    H h197(clk,reset,4'h1,2176'h0,h3InCommitment[197],Hstart[197],restart[197],groupNum,hashValue[197],en_end[197]);
    H h198(clk,reset,4'h1,2176'h0,h3InCommitment[198],Hstart[198],restart[198],groupNum,hashValue[198],en_end[198]);
    H h199(clk,reset,4'h1,2176'h0,h3InCommitment[199],Hstart[199],restart[199],groupNum,hashValue[199],en_end[199]);
    H h200(clk,reset,4'h1,2176'h0,h3InCommitment[200],Hstart[200],restart[200],groupNum,hashValue[200],en_end[200]);
    H h201(clk,reset,4'h1,2176'h0,h3InCommitment[201],Hstart[201],restart[201],groupNum,hashValue[201],en_end[201]);
    H h202(clk,reset,4'h1,2176'h0,h3InCommitment[202],Hstart[202],restart[202],groupNum,hashValue[202],en_end[202]);
    H h203(clk,reset,4'h1,2176'h0,h3InCommitment[203],Hstart[203],restart[203],groupNum,hashValue[203],en_end[203]);
    H h204(clk,reset,4'h1,2176'h0,h3InCommitment[204],Hstart[204],restart[204],groupNum,hashValue[204],en_end[204]);
    H h205(clk,reset,4'h1,2176'h0,h3InCommitment[205],Hstart[205],restart[205],groupNum,hashValue[205],en_end[205]);
    H h206(clk,reset,4'h1,2176'h0,h3InCommitment[206],Hstart[206],restart[206],groupNum,hashValue[206],en_end[206]);
    H h207(clk,reset,4'h1,2176'h0,h3InCommitment[207],Hstart[207],restart[207],groupNum,hashValue[207],en_end[207]);
    H h208(clk,reset,4'h1,2176'h0,h3InCommitment[208],Hstart[208],restart[208],groupNum,hashValue[208],en_end[208]);
    H h209(clk,reset,4'h1,2176'h0,h3InCommitment[209],Hstart[209],restart[209],groupNum,hashValue[209],en_end[209]);
    H h210(clk,reset,4'h1,2176'h0,h3InCommitment[210],Hstart[210],restart[210],groupNum,hashValue[210],en_end[210]);
    H h211(clk,reset,4'h1,2176'h0,h3InCommitment[211],Hstart[211],restart[211],groupNum,hashValue[211],en_end[211]);
    H h212(clk,reset,4'h1,2176'h0,h3InCommitment[212],Hstart[212],restart[212],groupNum,hashValue[212],en_end[212]);
    H h213(clk,reset,4'h1,2176'h0,h3InCommitment[213],Hstart[213],restart[213],groupNum,hashValue[213],en_end[213]);
    H h214(clk,reset,4'h1,2176'h0,h3InCommitment[214],Hstart[214],restart[214],groupNum,hashValue[214],en_end[214]);
    H h215(clk,reset,4'h1,2176'h0,h3InCommitment[215],Hstart[215],restart[215],groupNum,hashValue[215],en_end[215]);
    H h216(clk,reset,4'h1,2176'h0,h3InCommitment[216],Hstart[216],restart[216],groupNum,hashValue[216],en_end[216]);
    H h217(clk,reset,4'h1,2176'h0,h3InCommitment[217],Hstart[217],restart[217],groupNum,hashValue[217],en_end[217]);
    H h218(clk,reset,4'h1,2176'h0,h3InCommitment[218],Hstart[218],restart[218],groupNum,hashValue[218],en_end[218]);
    H h219(clk,reset,4'h1,2176'h0,h3InCommitment[219],Hstart[219],restart[219],groupNum,hashValue[219],en_end[219]);
    H h220(clk,reset,4'h1,2176'h0,h3InCommitment[220],Hstart[220],restart[220],groupNum,hashValue[220],en_end[220]);
    H h221(clk,reset,4'h1,2176'h0,h3InCommitment[221],Hstart[221],restart[221],groupNum,hashValue[221],en_end[221]);
    H h222(clk,reset,4'h1,2176'h0,h3InCommitment[222],Hstart[222],restart[222],groupNum,hashValue[222],en_end[222]);
    H h223(clk,reset,4'h1,2176'h0,h3InCommitment[223],Hstart[223],restart[223],groupNum,hashValue[223],en_end[223]);
    H h224(clk,reset,4'h1,2176'h0,h3InCommitment[224],Hstart[224],restart[224],groupNum,hashValue[224],en_end[224]);
    H h225(clk,reset,4'h1,2176'h0,h3InCommitment[225],Hstart[225],restart[225],groupNum,hashValue[225],en_end[225]);
    H h226(clk,reset,4'h1,2176'h0,h3InCommitment[226],Hstart[226],restart[226],groupNum,hashValue[226],en_end[226]);
    H h227(clk,reset,4'h1,2176'h0,h3InCommitment[227],Hstart[227],restart[227],groupNum,hashValue[227],en_end[227]);
    H h228(clk,reset,4'h1,2176'h0,h3InCommitment[228],Hstart[228],restart[228],groupNum,hashValue[228],en_end[228]);
    H h229(clk,reset,4'h1,2176'h0,h3InCommitment[229],Hstart[229],restart[229],groupNum,hashValue[229],en_end[229]);
    H h230(clk,reset,4'h1,2176'h0,h3InCommitment[230],Hstart[230],restart[230],groupNum,hashValue[230],en_end[230]);
    H h231(clk,reset,4'h1,2176'h0,h3InCommitment[231],Hstart[231],restart[231],groupNum,hashValue[231],en_end[231]);
    H h232(clk,reset,4'h1,2176'h0,h3InCommitment[232],Hstart[232],restart[232],groupNum,hashValue[232],en_end[232]);
    H h233(clk,reset,4'h1,2176'h0,h3InCommitment[233],Hstart[233],restart[233],groupNum,hashValue[233],en_end[233]);
    H h234(clk,reset,4'h1,2176'h0,h3InCommitment[234],Hstart[234],restart[234],groupNum,hashValue[234],en_end[234]);
    H h235(clk,reset,4'h1,2176'h0,h3InCommitment[235],Hstart[235],restart[235],groupNum,hashValue[235],en_end[235]);
    H h236(clk,reset,4'h1,2176'h0,h3InCommitment[236],Hstart[236],restart[236],groupNum,hashValue[236],en_end[236]);
    H h237(clk,reset,4'h1,2176'h0,h3InCommitment[237],Hstart[237],restart[237],groupNum,hashValue[237],en_end[237]);
    H h238(clk,reset,4'h1,2176'h0,h3InCommitment[238],Hstart[238],restart[238],groupNum,hashValue[238],en_end[238]);
    H h239(clk,reset,4'h1,2176'h0,h3InCommitment[239],Hstart[239],restart[239],groupNum,hashValue[239],en_end[239]);
    H h240(clk,reset,4'h1,2176'h0,h3InCommitment[240],Hstart[240],restart[240],groupNum,hashValue[240],en_end[240]);
    H h241(clk,reset,4'h1,2176'h0,h3InCommitment[241],Hstart[241],restart[241],groupNum,hashValue[241],en_end[241]);
    H h242(clk,reset,4'h1,2176'h0,h3InCommitment[242],Hstart[242],restart[242],groupNum,hashValue[242],en_end[242]);
    H h243(clk,reset,4'h1,2176'h0,h3InCommitment[243],Hstart[243],restart[243],groupNum,hashValue[243],en_end[243]);
    H h244(clk,reset,4'h1,2176'h0,h3InCommitment[244],Hstart[244],restart[244],groupNum,hashValue[244],en_end[244]);
    H h245(clk,reset,4'h1,2176'h0,h3InCommitment[245],Hstart[245],restart[245],groupNum,hashValue[245],en_end[245]);
    H h246(clk,reset,4'h1,2176'h0,h3InCommitment[246],Hstart[246],restart[246],groupNum,hashValue[246],en_end[246]);
    H h247(clk,reset,4'h1,2176'h0,h3InCommitment[247],Hstart[247],restart[247],groupNum,hashValue[247],en_end[247]);
    H h248(clk,reset,4'h1,2176'h0,h3InCommitment[248],Hstart[248],restart[248],groupNum,hashValue[248],en_end[248]);
    H h249(clk,reset,4'h1,2176'h0,h3InCommitment[249],Hstart[249],restart[249],groupNum,hashValue[249],en_end[249]);
    H h250(clk,reset,4'h1,2176'h0,h3InCommitment[250],Hstart[250],restart[250],groupNum,hashValue[250],en_end[250]);
    H h251(clk,reset,4'h1,2176'h0,h3InCommitment[251],Hstart[251],restart[251],groupNum,hashValue[251],en_end[251]);
    H h252(clk,reset,4'h1,2176'h0,h3InCommitment[252],Hstart[252],restart[252],groupNum,hashValue[252],en_end[252]);
    H h253(clk,reset,4'h1,2176'h0,h3InCommitment[253],Hstart[253],restart[253],groupNum,hashValue[253],en_end[253]);
    H h254(clk,reset,4'h1,2176'h0,h3InCommitment[254],Hstart[254],restart[254],groupNum,hashValue[254],en_end[254]);
    H h255(clk,reset,4'h1,2176'h0,h3InCommitment[255],Hstart[255],restart[255],groupNum,hashValue[255],en_end[255]);
    H h256(clk,reset,4'h1,2176'h0,h3InCommitment[256],Hstart[256],restart[256],groupNum,hashValue[256],en_end[256]);
    H h257(clk,reset,4'h1,2176'h0,h3InCommitment[257],Hstart[257],restart[257],groupNum,hashValue[257],en_end[257]);
    H h258(clk,reset,4'h1,2176'h0,h3InCommitment[258],Hstart[258],restart[258],groupNum,hashValue[258],en_end[258]);
    H h259(clk,reset,4'h1,2176'h0,h3InCommitment[259],Hstart[259],restart[259],groupNum,hashValue[259],en_end[259]);
    H h260(clk,reset,4'h1,2176'h0,h3InCommitment[260],Hstart[260],restart[260],groupNum,hashValue[260],en_end[260]);
    H h261(clk,reset,4'h1,2176'h0,h3InCommitment[261],Hstart[261],restart[261],groupNum,hashValue[261],en_end[261]);
    H h262(clk,reset,4'h1,2176'h0,h3InCommitment[262],Hstart[262],restart[262],groupNum,hashValue[262],en_end[262]);
    H h263(clk,reset,4'h1,2176'h0,h3InCommitment[263],Hstart[263],restart[263],groupNum,hashValue[263],en_end[263]);
    H h264(clk,reset,4'h1,2176'h0,h3InCommitment[264],Hstart[264],restart[264],groupNum,hashValue[264],en_end[264]);
    H h265(clk,reset,4'h1,2176'h0,h3InCommitment[265],Hstart[265],restart[265],groupNum,hashValue[265],en_end[265]);
    H h266(clk,reset,4'h1,2176'h0,h3InCommitment[266],Hstart[266],restart[266],groupNum,hashValue[266],en_end[266]);
    H h267(clk,reset,4'h1,2176'h0,h3InCommitment[267],Hstart[267],restart[267],groupNum,hashValue[267],en_end[267]);
    H h268(clk,reset,4'h1,2176'h0,h3InCommitment[268],Hstart[268],restart[268],groupNum,hashValue[268],en_end[268]);
    H h269(clk,reset,4'h1,2176'h0,h3InCommitment[269],Hstart[269],restart[269],groupNum,hashValue[269],en_end[269]);
    H h270(clk,reset,4'h1,2176'h0,h3InCommitment[270],Hstart[270],restart[270],groupNum,hashValue[270],en_end[270]);
    H h271(clk,reset,4'h1,2176'h0,h3InCommitment[271],Hstart[271],restart[271],groupNum,hashValue[271],en_end[271]);
    H h272(clk,reset,4'h1,2176'h0,h3InCommitment[272],Hstart[272],restart[272],groupNum,hashValue[272],en_end[272]);
    H h273(clk,reset,4'h1,2176'h0,h3InCommitment[273],Hstart[273],restart[273],groupNum,hashValue[273],en_end[273]);
    H h274(clk,reset,4'h1,2176'h0,h3InCommitment[274],Hstart[274],restart[274],groupNum,hashValue[274],en_end[274]);
    H h275(clk,reset,4'h1,2176'h0,h3InCommitment[275],Hstart[275],restart[275],groupNum,hashValue[275],en_end[275]);
    H h276(clk,reset,4'h1,2176'h0,h3InCommitment[276],Hstart[276],restart[276],groupNum,hashValue[276],en_end[276]);
    H h277(clk,reset,4'h1,2176'h0,h3InCommitment[277],Hstart[277],restart[277],groupNum,hashValue[277],en_end[277]);
    H h278(clk,reset,4'h1,2176'h0,h3InCommitment[278],Hstart[278],restart[278],groupNum,hashValue[278],en_end[278]);
    H h279(clk,reset,4'h1,2176'h0,h3InCommitment[279],Hstart[279],restart[279],groupNum,hashValue[279],en_end[279]);
    H h280(clk,reset,4'h1,2176'h0,h3InCommitment[280],Hstart[280],restart[280],groupNum,hashValue[280],en_end[280]);
    H h281(clk,reset,4'h1,2176'h0,h3InCommitment[281],Hstart[281],restart[281],groupNum,hashValue[281],en_end[281]);
    H h282(clk,reset,4'h1,2176'h0,h3InCommitment[282],Hstart[282],restart[282],groupNum,hashValue[282],en_end[282]);
    H h283(clk,reset,4'h1,2176'h0,h3InCommitment[283],Hstart[283],restart[283],groupNum,hashValue[283],en_end[283]);
    H h284(clk,reset,4'h1,2176'h0,h3InCommitment[284],Hstart[284],restart[284],groupNum,hashValue[284],en_end[284]);
    H h285(clk,reset,4'h1,2176'h0,h3InCommitment[285],Hstart[285],restart[285],groupNum,hashValue[285],en_end[285]);
    H h286(clk,reset,4'h1,2176'h0,h3InCommitment[286],Hstart[286],restart[286],groupNum,hashValue[286],en_end[286]);
    H h287(clk,reset,4'h1,2176'h0,h3InCommitment[287],Hstart[287],restart[287],groupNum,hashValue[287],en_end[287]);
    H h288(clk,reset,4'h1,2176'h0,h3InCommitment[288],Hstart[288],restart[288],groupNum,hashValue[288],en_end[288]);
    H h289(clk,reset,4'h1,2176'h0,h3InCommitment[289],Hstart[289],restart[289],groupNum,hashValue[289],en_end[289]);
    H h290(clk,reset,4'h1,2176'h0,h3InCommitment[290],Hstart[290],restart[290],groupNum,hashValue[290],en_end[290]);
    H h291(clk,reset,4'h1,2176'h0,h3InCommitment[291],Hstart[291],restart[291],groupNum,hashValue[291],en_end[291]);
    H h292(clk,reset,4'h1,2176'h0,h3InCommitment[292],Hstart[292],restart[292],groupNum,hashValue[292],en_end[292]);
    H h293(clk,reset,4'h1,2176'h0,h3InCommitment[293],Hstart[293],restart[293],groupNum,hashValue[293],en_end[293]);
    H h294(clk,reset,4'h1,2176'h0,h3InCommitment[294],Hstart[294],restart[294],groupNum,hashValue[294],en_end[294]);
    H h295(clk,reset,4'h1,2176'h0,h3InCommitment[295],Hstart[295],restart[295],groupNum,hashValue[295],en_end[295]);
    H h296(clk,reset,4'h1,2176'h0,h3InCommitment[296],Hstart[296],restart[296],groupNum,hashValue[296],en_end[296]);
    H h297(clk,reset,4'h1,2176'h0,h3InCommitment[297],Hstart[297],restart[297],groupNum,hashValue[297],en_end[297]);
    H h298(clk,reset,4'h1,2176'h0,h3InCommitment[298],Hstart[298],restart[298],groupNum,hashValue[298],en_end[298]);
    H h299(clk,reset,4'h1,2176'h0,h3InCommitment[299],Hstart[299],restart[299],groupNum,hashValue[299],en_end[299]);
    H h300(clk,reset,4'h1,2176'h0,h3InCommitment[300],Hstart[300],restart[300],groupNum,hashValue[300],en_end[300]);
endmodule