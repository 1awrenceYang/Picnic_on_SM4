`timescale 1ns / 1ps
module CalculateT_result(
    input [7:0] a,
    output [7:0] final
    );
    
wire T_result0, T_result1, T_result2, T_result3, T_result4;
wire T_result10, T_result11, T_result12, T_result13, T_result14;
wire T_result20, T_result21, T_result22, T_result23, T_result24;
wire T_result30, T_result31, T_result32, T_result33, T_result34;
wire T_result40, T_result41, T_result42, T_result43, T_result44;
wire T_result50, T_result51, T_result52, T_result53, T_result54;
wire T_result60, T_result61, T_result62, T_result63, T_result64;
wire T_result70, T_result71, T_result72, T_result73, T_result74;

assign T_result0= (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]) ^ (a[4]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[3]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]);
assign T_result1=(a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]);
assign T_result2=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]);
assign T_result3=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]);
assign T_result4=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign T_result10=(a[7]) ^ (a[6]) ^ (a[7]) ^ (a[6]&a[7]) ^ (a[5]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]) ^ (a[4]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]);
assign T_result11=(a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]);
assign T_result12=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]);
assign T_result13=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]);
assign T_result14=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign T_result20=(a[6]) ^ (a[5]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]);
assign T_result21=(a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]);
assign T_result22=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]);
assign T_result23=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]);
assign T_result24=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign T_result30=(a[6]) ^ (a[6]) ^ (a[7]) ^ (a[6]&a[7]) ^ (a[5]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]);
assign T_result31=(a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[0]) ^ (a[7]) ^ (a[0]&a[7]);
assign T_result32=(a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]);
assign T_result33=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]);
assign T_result34=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign T_result40=(a[6]) ^ (a[5]) ^ (a[5]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[3]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[2]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]);
assign T_result41=(a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]);
assign T_result42=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]);
assign T_result43=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]&a[7]);
assign T_result44=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]);

assign T_result50=(a[7]) ^ (a[6]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[3]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]);
assign T_result51=(a[1]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]);
assign T_result52=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]);
assign T_result53=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]);
assign T_result54=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign T_result60=(a[7]) ^ (a[6]) ^ (a[5]) ^ (a[5]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[5]) ^ (a[6]) ^ (a[5]&a[6]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[4]) ^ (a[5]) ^ (a[4]&a[5]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]);
assign T_result61=(a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]);
assign T_result62=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]);
assign T_result63=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]);
assign T_result64=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign T_result70=(a[6]) ^ (a[6]) ^ (a[7]) ^ (a[6]&a[7]) ^ (a[5]) ^ (a[7]) ^ (a[5]&a[7]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[4]) ^ (a[6]) ^ (a[4]&a[6]) ^ (a[7]) ^ (a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[3]) ^ (a[3]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[3]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[3]) ^ (a[4]) ^ (a[3]&a[4]) ^ (a[5]) ^ (a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[2]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[2]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]);
assign T_result71=(a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]) ^ (a[3]) ^ (a[2]&a[3]) ^ (a[4]) ^ (a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[1]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[1]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]);
assign T_result72=(a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]) ^ (a[2]) ^ (a[1]&a[2]) ^ (a[3]) ^ (a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[0]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[0]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]);
assign T_result73=(a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[2]&a[4]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[2]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]);
assign T_result74=(a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[4]&a[6]&a[7]) ^ (a[0]&a[4]&a[6]&a[7]) ^ (a[1]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[6]&a[7]) ^ (a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]&a[7]) ^ (a[5]&a[6]&a[7]) ^ (a[0]&a[5]&a[6]&a[7]) ^ (a[1]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[5]&a[6]&a[7]) ^ (a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]&a[7]) ^ (a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]&a[7]) ^ (a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[6]&a[7]) ^ (a[0]&a[6]&a[7]) ^ (a[1]&a[6]&a[7]) ^ (a[0]&a[1]&a[6]&a[7]) ^ (a[2]&a[6]&a[7]) ^ (a[0]&a[2]&a[6]&a[7]) ^ (a[1]&a[2]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[6]&a[7]) ^ (a[3]&a[6]&a[7]) ^ (a[0]&a[3]&a[6]&a[7]) ^ (a[1]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[3]&a[6]&a[7]) ^ (a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[2]&a[3]&a[6]&a[7]) ^ (a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[7]) ^ (a[0]&a[7]) ^ (a[1]&a[7]) ^ (a[0]&a[1]&a[7]) ^ (a[2]&a[7]) ^ (a[0]&a[2]&a[7]) ^ (a[1]&a[2]&a[7]) ^ (a[0]&a[1]&a[2]&a[7]) ^ (a[3]&a[7]) ^ (a[0]&a[3]&a[7]) ^ (a[1]&a[3]&a[7]) ^ (a[0]&a[1]&a[3]&a[7]) ^ (a[2]&a[3]&a[7]) ^ (a[0]&a[2]&a[3]&a[7]) ^ (a[1]&a[2]&a[3]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[7]) ^ (a[4]&a[7]) ^ (a[0]&a[4]&a[7]) ^ (a[1]&a[4]&a[7]) ^ (a[0]&a[1]&a[4]&a[7]) ^ (a[2]&a[4]&a[7]) ^ (a[0]&a[2]&a[4]&a[7]) ^ (a[1]&a[2]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[7]) ^ (a[3]&a[4]&a[7]) ^ (a[0]&a[3]&a[4]&a[7]) ^ (a[1]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[7]) ^ (a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[7]) ^ (a[5]&a[7]) ^ (a[0]&a[5]&a[7]) ^ (a[1]&a[5]&a[7]) ^ (a[0]&a[1]&a[5]&a[7]) ^ (a[2]&a[5]&a[7]) ^ (a[0]&a[2]&a[5]&a[7]) ^ (a[1]&a[2]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[5]&a[7]) ^ (a[3]&a[5]&a[7]) ^ (a[0]&a[3]&a[5]&a[7]) ^ (a[1]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[5]&a[7]) ^ (a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[7]) ^ (a[4]&a[5]&a[7]) ^ (a[0]&a[4]&a[5]&a[7]) ^ (a[1]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[4]&a[5]&a[7]) ^ (a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[7]) ^ (a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[7]) ^ (a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[7]) ^ (a[0]) ^ (a[1]) ^ (a[0]&a[1]) ^ (a[2]) ^ (a[0]&a[2]) ^ (a[1]&a[2]) ^ (a[0]&a[1]&a[2]) ^ (a[3]) ^ (a[0]&a[3]) ^ (a[1]&a[3]) ^ (a[0]&a[1]&a[3]) ^ (a[2]&a[3]) ^ (a[0]&a[2]&a[3]) ^ (a[1]&a[2]&a[3]) ^ (a[0]&a[1]&a[2]&a[3]) ^ (a[4]) ^ (a[0]&a[4]) ^ (a[1]&a[4]) ^ (a[0]&a[1]&a[4]) ^ (a[2]&a[4]) ^ (a[0]&a[2]&a[4]) ^ (a[1]&a[2]&a[4]) ^ (a[0]&a[1]&a[2]&a[4]) ^ (a[3]&a[4]) ^ (a[0]&a[3]&a[4]) ^ (a[1]&a[3]&a[4]) ^ (a[0]&a[1]&a[3]&a[4]) ^ (a[2]&a[3]&a[4]) ^ (a[0]&a[2]&a[3]&a[4]) ^ (a[1]&a[2]&a[3]&a[4]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]) ^ (a[5]) ^ (a[0]&a[5]) ^ (a[1]&a[5]) ^ (a[0]&a[1]&a[5]) ^ (a[2]&a[5]) ^ (a[0]&a[2]&a[5]) ^ (a[1]&a[2]&a[5]) ^ (a[0]&a[1]&a[2]&a[5]) ^ (a[3]&a[5]) ^ (a[0]&a[3]&a[5]) ^ (a[1]&a[3]&a[5]) ^ (a[0]&a[1]&a[3]&a[5]) ^ (a[2]&a[3]&a[5]) ^ (a[0]&a[2]&a[3]&a[5]) ^ (a[1]&a[2]&a[3]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]) ^ (a[4]&a[5]) ^ (a[0]&a[4]&a[5]) ^ (a[1]&a[4]&a[5]) ^ (a[0]&a[1]&a[4]&a[5]) ^ (a[2]&a[4]&a[5]) ^ (a[0]&a[2]&a[4]&a[5]) ^ (a[1]&a[2]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]) ^ (a[3]&a[4]&a[5]) ^ (a[0]&a[3]&a[4]&a[5]) ^ (a[1]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]) ^ (a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]) ^ (a[6]) ^ (a[0]&a[6]) ^ (a[1]&a[6]) ^ (a[0]&a[1]&a[6]) ^ (a[2]&a[6]) ^ (a[0]&a[2]&a[6]) ^ (a[1]&a[2]&a[6]) ^ (a[0]&a[1]&a[2]&a[6]) ^ (a[3]&a[6]) ^ (a[0]&a[3]&a[6]) ^ (a[1]&a[3]&a[6]) ^ (a[0]&a[1]&a[3]&a[6]) ^ (a[2]&a[3]&a[6]) ^ (a[0]&a[2]&a[3]&a[6]) ^ (a[1]&a[2]&a[3]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[6]) ^ (a[4]&a[6]) ^ (a[0]&a[4]&a[6]) ^ (a[1]&a[4]&a[6]) ^ (a[0]&a[1]&a[4]&a[6]) ^ (a[2]&a[4]&a[6]) ^ (a[0]&a[2]&a[4]&a[6]) ^ (a[1]&a[2]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[6]) ^ (a[3]&a[4]&a[6]) ^ (a[0]&a[3]&a[4]&a[6]) ^ (a[1]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[6]) ^ (a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[6]) ^ (a[5]&a[6]) ^ (a[0]&a[5]&a[6]) ^ (a[1]&a[5]&a[6]) ^ (a[0]&a[1]&a[5]&a[6]) ^ (a[2]&a[5]&a[6]) ^ (a[0]&a[2]&a[5]&a[6]) ^ (a[1]&a[2]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[5]&a[6]) ^ (a[3]&a[5]&a[6]) ^ (a[0]&a[3]&a[5]&a[6]) ^ (a[1]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[5]&a[6]) ^ (a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[5]&a[6]) ^ (a[4]&a[5]&a[6]) ^ (a[0]&a[4]&a[5]&a[6]) ^ (a[1]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[4]&a[5]&a[6]) ^ (a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[4]&a[5]&a[6]) ^ (a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[3]&a[4]&a[5]&a[6]) ^ (a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[1]&a[2]&a[3]&a[4]&a[5]&a[6]) ^ (a[0]&a[1]&a[2]&a[3]&a[4]&a[5]&a[6]);

assign final[0]=T_result0^T_result1^T_result2^T_result3^T_result4;
assign final[1]=T_result10^T_result11^T_result12^T_result13^T_result14;
assign final[2]=T_result20^T_result21^T_result22^T_result23^T_result24;
assign final[3]=T_result30^T_result31^T_result32^T_result33^T_result34;
assign final[4]=T_result40^T_result41^T_result42^T_result43^T_result44;
assign final[5]=T_result50^T_result51^T_result52^T_result53^T_result54;
assign final[6]=T_result60^T_result61^T_result62^T_result63^T_result64;
assign final[7]=T_result70^T_result71^T_result72^T_result73^T_result74;
endmodule

module Compute_lambda_I(
    input [7:0] masked_input,
    output [254:0] Lambda_I
);
    
assign Lambda_I[0]=masked_input[0];
assign Lambda_I[1]=masked_input[1];
assign Lambda_I[2]=masked_input[1] & masked_input[0];
assign Lambda_I[3]=masked_input[2];
assign Lambda_I[4]=masked_input[2] & masked_input[0];
assign Lambda_I[5]=masked_input[2] & masked_input[1];
assign Lambda_I[6]=masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[7]=masked_input[3];
assign Lambda_I[8]=masked_input[3] & masked_input[0];
assign Lambda_I[9]=masked_input[3] & masked_input[1];
assign Lambda_I[10]=masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[11]=masked_input[3] & masked_input[2];
assign Lambda_I[12]=masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[13]=masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[14]=masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[15]=masked_input[4];
assign Lambda_I[16]=masked_input[4] & masked_input[0];
assign Lambda_I[17]=masked_input[4] & masked_input[1];
assign Lambda_I[18]=masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[19]=masked_input[4] & masked_input[2];
assign Lambda_I[20]=masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[21]=masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[22]=masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[23]=masked_input[4] & masked_input[3];
assign Lambda_I[24]=masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[25]=masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[26]=masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[27]=masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[28]=masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[29]=masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[30]=masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[31]=masked_input[5];
assign Lambda_I[32]=masked_input[5] & masked_input[0];
assign Lambda_I[33]=masked_input[5] & masked_input[1];
assign Lambda_I[34]=masked_input[5] & masked_input[1] & masked_input[0];
assign Lambda_I[35]=masked_input[5] & masked_input[2];
assign Lambda_I[36]=masked_input[5] & masked_input[2] & masked_input[0];
assign Lambda_I[37]=masked_input[5] & masked_input[2] & masked_input[1];
assign Lambda_I[38]=masked_input[5] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[39]=masked_input[5] & masked_input[3];
assign Lambda_I[40]=masked_input[5] & masked_input[3] & masked_input[0];
assign Lambda_I[41]=masked_input[5] & masked_input[3] & masked_input[1];
assign Lambda_I[42]=masked_input[5] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[43]=masked_input[5] & masked_input[3] & masked_input[2];
assign Lambda_I[44]=masked_input[5] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[45]=masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[46]=masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[47]=masked_input[5] & masked_input[4];
assign Lambda_I[48]=masked_input[5] & masked_input[4] & masked_input[0];
assign Lambda_I[49]=masked_input[5] & masked_input[4] & masked_input[1];
assign Lambda_I[50]=masked_input[5] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[51]=masked_input[5] & masked_input[4] & masked_input[2];
assign Lambda_I[52]=masked_input[5] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[53]=masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[54]=masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[55]=masked_input[5] & masked_input[4] & masked_input[3];
assign Lambda_I[56]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[57]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[58]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[59]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[60]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[61]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[62]=masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[63]=masked_input[6];
assign Lambda_I[64]=masked_input[6] & masked_input[0];
assign Lambda_I[65]=masked_input[6] & masked_input[1];
assign Lambda_I[66]=masked_input[6] & masked_input[1] & masked_input[0];
assign Lambda_I[67]=masked_input[6] & masked_input[2];
assign Lambda_I[68]=masked_input[6] & masked_input[2] & masked_input[0];
assign Lambda_I[69]=masked_input[6] & masked_input[2] & masked_input[1];
assign Lambda_I[70]=masked_input[6] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[71]=masked_input[6] & masked_input[3];
assign Lambda_I[72]=masked_input[6] & masked_input[3] & masked_input[0];
assign Lambda_I[73]=masked_input[6] & masked_input[3] & masked_input[1];
assign Lambda_I[74]=masked_input[6] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[75]=masked_input[6] & masked_input[3] & masked_input[2];
assign Lambda_I[76]=masked_input[6] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[77]=masked_input[6] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[78]=masked_input[6] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[79]=masked_input[6] & masked_input[4];
assign Lambda_I[80]=masked_input[6] & masked_input[4] & masked_input[0];
assign Lambda_I[81]=masked_input[6] & masked_input[4] & masked_input[1];
assign Lambda_I[82]=masked_input[6] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[83]=masked_input[6] & masked_input[4] & masked_input[2];
assign Lambda_I[84]=masked_input[6] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[85]=masked_input[6] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[86]=masked_input[6] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[87]=masked_input[6] & masked_input[4] & masked_input[3];
assign Lambda_I[88]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[89]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[90]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[91]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[92]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[93]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[94]=masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[95]=masked_input[6] & masked_input[5];
assign Lambda_I[96]=masked_input[6] & masked_input[5] & masked_input[0];
assign Lambda_I[97]=masked_input[6] & masked_input[5] & masked_input[1];
assign Lambda_I[98]=masked_input[6] & masked_input[5] & masked_input[1] & masked_input[0];
assign Lambda_I[99]=masked_input[6] & masked_input[5] & masked_input[2];
assign Lambda_I[100]=masked_input[6] & masked_input[5] & masked_input[2] & masked_input[0];
assign Lambda_I[101]=masked_input[6] & masked_input[5] & masked_input[2] & masked_input[1];
assign Lambda_I[102]=masked_input[6] & masked_input[5] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[103]=masked_input[6] & masked_input[5] & masked_input[3];
assign Lambda_I[104]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[0];
assign Lambda_I[105]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[1];
assign Lambda_I[106]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[107]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2];
assign Lambda_I[108]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[109]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[110]=masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[111]=masked_input[6] & masked_input[5] & masked_input[4];
assign Lambda_I[112]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[0];
assign Lambda_I[113]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[1];
assign Lambda_I[114]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[115]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2];
assign Lambda_I[116]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[117]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[118]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[119]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3];
assign Lambda_I[120]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[121]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[122]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[123]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[124]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[125]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[126]=masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[127]=masked_input[7];
assign Lambda_I[128]=masked_input[7] & masked_input[0];
assign Lambda_I[129]=masked_input[7] & masked_input[1];
assign Lambda_I[130]=masked_input[7] & masked_input[1] & masked_input[0];
assign Lambda_I[131]=masked_input[7] & masked_input[2];
assign Lambda_I[132]=masked_input[7] & masked_input[2] & masked_input[0];
assign Lambda_I[133]=masked_input[7] & masked_input[2] & masked_input[1];
assign Lambda_I[134]=masked_input[7] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[135]=masked_input[7] & masked_input[3];
assign Lambda_I[136]=masked_input[7] & masked_input[3] & masked_input[0];
assign Lambda_I[137]=masked_input[7] & masked_input[3] & masked_input[1];
assign Lambda_I[138]=masked_input[7] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[139]=masked_input[7] & masked_input[3] & masked_input[2];
assign Lambda_I[140]=masked_input[7] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[141]=masked_input[7] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[142]=masked_input[7] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[143]=masked_input[7] & masked_input[4];
assign Lambda_I[144]=masked_input[7] & masked_input[4] & masked_input[0];
assign Lambda_I[145]=masked_input[7] & masked_input[4] & masked_input[1];
assign Lambda_I[146]=masked_input[7] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[147]=masked_input[7] & masked_input[4] & masked_input[2];
assign Lambda_I[148]=masked_input[7] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[149]=masked_input[7] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[150]=masked_input[7] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[151]=masked_input[7] & masked_input[4] & masked_input[3];
assign Lambda_I[152]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[153]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[154]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[155]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[156]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[157]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[158]=masked_input[7] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[159]=masked_input[7] & masked_input[5];
assign Lambda_I[160]=masked_input[7] & masked_input[5] & masked_input[0];
assign Lambda_I[161]=masked_input[7] & masked_input[5] & masked_input[1];
assign Lambda_I[162]=masked_input[7] & masked_input[5] & masked_input[1] & masked_input[0];
assign Lambda_I[163]=masked_input[7] & masked_input[5] & masked_input[2];
assign Lambda_I[164]=masked_input[7] & masked_input[5] & masked_input[2] & masked_input[0];
assign Lambda_I[165]=masked_input[7] & masked_input[5] & masked_input[2] & masked_input[1];
assign Lambda_I[166]=masked_input[7] & masked_input[5] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[167]=masked_input[7] & masked_input[5] & masked_input[3];
assign Lambda_I[168]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[0];
assign Lambda_I[169]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[1];
assign Lambda_I[170]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[171]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[2];
assign Lambda_I[172]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[173]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[174]=masked_input[7] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[175]=masked_input[7] & masked_input[5] & masked_input[4];
assign Lambda_I[176]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[0];
assign Lambda_I[177]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[1];
assign Lambda_I[178]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[179]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[2];
assign Lambda_I[180]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[181]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[182]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[183]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3];
assign Lambda_I[184]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[185]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[186]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[187]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[188]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[189]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[190]=masked_input[7] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[191]=masked_input[7] & masked_input[6];
assign Lambda_I[192]=masked_input[7] & masked_input[6] & masked_input[0];
assign Lambda_I[193]=masked_input[7] & masked_input[6] & masked_input[1];
assign Lambda_I[194]=masked_input[7] & masked_input[6] & masked_input[1] & masked_input[0];
assign Lambda_I[195]=masked_input[7] & masked_input[6] & masked_input[2];
assign Lambda_I[196]=masked_input[7] & masked_input[6] & masked_input[2] & masked_input[0];
assign Lambda_I[197]=masked_input[7] & masked_input[6] & masked_input[2] & masked_input[1];
assign Lambda_I[198]=masked_input[7] & masked_input[6] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[199]=masked_input[7] & masked_input[6] & masked_input[3];
assign Lambda_I[200]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[0];
assign Lambda_I[201]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[1];
assign Lambda_I[202]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[203]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[2];
assign Lambda_I[204]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[205]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[206]=masked_input[7] & masked_input[6] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[207]=masked_input[7] & masked_input[6] & masked_input[4];
assign Lambda_I[208]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[0];
assign Lambda_I[209]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[1];
assign Lambda_I[210]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[211]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[2];
assign Lambda_I[212]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[213]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[214]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[215]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3];
assign Lambda_I[216]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[217]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[218]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[219]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[220]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[221]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[222]=masked_input[7] & masked_input[6] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[223]=masked_input[7] & masked_input[6] & masked_input[5];
assign Lambda_I[224]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[0];
assign Lambda_I[225]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[1];
assign Lambda_I[226]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[1] & masked_input[0];
assign Lambda_I[227]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[2];
assign Lambda_I[228]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[2] & masked_input[0];
assign Lambda_I[229]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[2] & masked_input[1];
assign Lambda_I[230]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[231]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3];
assign Lambda_I[232]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[0];
assign Lambda_I[233]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[1];
assign Lambda_I[234]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[235]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2];
assign Lambda_I[236]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[237]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[238]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[239]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4];
assign Lambda_I[240]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[0];
assign Lambda_I[241]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[1];
assign Lambda_I[242]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[1] & masked_input[0];
assign Lambda_I[243]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2];
assign Lambda_I[244]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[0];
assign Lambda_I[245]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1];
assign Lambda_I[246]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[2] & masked_input[1] & masked_input[0];
assign Lambda_I[247]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3];
assign Lambda_I[248]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[0];
assign Lambda_I[249]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1];
assign Lambda_I[250]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[1] & masked_input[0];
assign Lambda_I[251]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2];
assign Lambda_I[252]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[0];
assign Lambda_I[253]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1];
assign Lambda_I[254]=masked_input[7] & masked_input[6] & masked_input[5] & masked_input[4] & masked_input[3] & masked_input[2] & masked_input[1] & masked_input[0];
    
    
endmodule

module compute_aux_bits(
    input [31:0] xored_round_key,
    output [255*4-1:0] out
);
    wire [254:0] Lambda_I1, Lambda_I2, Lambda_I3, Lambda_I4;
    
    
    Compute_lambda_I compute1(xored_round_key[7:0], out[254:0]);
    Compute_lambda_I compute2(xored_round_key[15:8], out[509:255]);
    Compute_lambda_I compute3(xored_round_key[23:16], out[764:510]);
    Compute_lambda_I compute4(xored_round_key[31:24], out[1019:765]);
    
endmodule

module compute_aux_read_tapes(
    input clk,
    input rst,
    input [4:0] round,
    input [1:0] k,
    input start,
    input [1:0] operating_mode,//from 00-11 for compute_aux_sign_first_right, compute_aux_sign_first_left, 
    output [254:0] xor_result,
    output [254:0] xor_result2,
    output reg stop
);
// original value: e8db9ae7a5a937278b60d5ca371b1481
//after L_matrix: 008e202eb5214106ffa2cb69226450d6
//mpc_output_reg<=128'h008e202eb5214106ffa2cb69226450d6;
reg [10:0] ReadAddress;
reg [254:0] tape0_result;
reg [254:0] tape1_result;
reg [3:0] state;
reg [3:0] counter;
reg read_en;
wire [527:0] temp;
wire [527:0] tapes_xor_result;
wire [10:0] ReadAddress_wire;
tapes random_tapes 
(
  .clka(clk),    // input wire clka
  .ena(1'b0),      // input wire ena
  .wea(1'b0),      // input wire [0 : 0] wea
  .addra(11'b0),  // input wire [10 : 0] addra
  .dina(528'b0),    // input wire [527 : 0] dina
  .clkb(clk),    // input wire clkb
  .enb(read_en),      // input wire enb
  .addrb(ReadAddress),  // input wire [10 : 0] addrb
  .doutb(tapes_xor_result)  // output wire [527 : 0] doutb
);

    Get_Read_Address GRA1(round, k, ReadAddress_wire);
    
    always@(posedge clk or negedge rst)
    begin
        if(!rst)
            begin
                ReadAddress<=11'b0;
                tape0_result<=255'b0;
                tape1_result<=255'b0;
                state<=4'b0;
                counter<=4'b0;
                read_en<=1'b0;
                stop<=1'b0;
            end
        else
            begin
                if(operating_mode==2'd0)
                    begin
                        if(state==4'd0)
                            begin
                                stop<=1'b0;
                                if(start)
                                    begin
                                        ReadAddress<=ReadAddress_wire;
                                        read_en<=1'b1;
                                        state=4'd1;
                                    end
                            end
                            
                        else if(state==4'd1)
                            begin
                                if(counter==4'd15)
                                    begin
                                        tape0_result<=tape0_result^tapes_xor_result[255:1];
                                        tape1_result<=tape1_result^tapes_xor_result[511:257];
                                        state<=4'd2;
                                        
                                    end
                                else
                                    begin
                                        tape0_result<=tape0_result^tapes_xor_result[255:1];
                                        tape1_result<=tape1_result^tapes_xor_result[511:257];
                                        counter<=counter+1;
                                        ReadAddress<=ReadAddress+128;
                                    end
                            end
                            
                        else if(state==4'd2)
                            begin
                                state<=4'd3;
                                stop<=1'b1;
                                read_en<=1'b0;
                            end
                            
                        else if(state==4'd3)
                            begin
                                state<=4'd0;
                                stop<=1'b1;
                            end
                    end
                    
                else if(operating_mode==2'b1)
                    begin
                        if(state==4'd0)
                            begin
                                stop<=1'b0;
                                if(start)
                                    begin
                                        ReadAddress<=ReadAddress_wire;
                                        read_en<=1'b1;
                                        state=4'd1;
                                    end
                            end
                            
                        else if(state==4'd1)
                            begin
                                if(counter==4'd15)
                                    begin
                                        tape0_result<=tape0_result^tapes_xor_result[511:257];
                                        state<=4'd2;
                                    end
                                else
                                    begin
                                        tape0_result<=tape0_result^tapes_xor_result[511:257];
                                        counter<=counter+1;
                                        ReadAddress<=ReadAddress+128;
                                    end
                            end
                            
                        else if(state==4'd2)
                            begin
                                state<=4'd3;
                                stop<=1'b1;
                                read_en<=1'b0;
                            end
                            
                        else if(state==4'd3)
                            begin
                                state<=4'd0;
                                stop<=1'b1;
                            end
                    end
            end
    end


assign xor_result=tape0_result;
assign xor_result2=tape1_result;
endmodule

module compute_aux_write_aux1(
    input clk,
    input rst,
    input [254:0] data_in,
    input start,
    input [4:0] round,
    
    output  stop,
    output  [511:0] out
    //output [4:0] state_out
);

reg [6:0] WriteAddress, ReadAddress;
reg rwControl, read_en, write_en;
reg [511:0] data;
reg [3:0] state;
reg stop_reg;
wire [511:0] data_out;

assign out=data_out;
//assign state_out=state;
assign stop=stop_reg;


aux_bits aux 
(
  .clka(clk),    // input wire clka
  .ena(write_en),      // input wire ena
  .wea(rwControl),      // input wire [0 : 0] wea
  .addra(WriteAddress),  // input wire [6 : 0] addra
  .dina(data),    // input wire [511 : 0] dina
  .clkb(clk),    // input wire clkb
  .enb(read_en),      // input wire enb
  .addrb(ReadAddress),  // input wire [6 : 0] addrb
  .doutb(data_out)  // output wire [511 : 0] doutb
);
    
    
always@(posedge clk or negedge rst)
begin
    if(!rst)
        begin
            data<=512'b0;
            write_en<=1'b0;
            read_en<=1'b0;
            rwControl<=1'b0;
            state<=4'b0000;
            ReadAddress<=7'b0;
            WriteAddress<=7'b0;
        end
    else
        if(state==4'b0000)
            begin
                stop_reg<=0;
                if(start)
                begin

                    data<={256'b0, data_in, 1'b0};
                    state<=4'b0001;
                    rwControl<=1'b1;
                    write_en<=1'b1;
                    read_en<=1'b0;

                case(round)
                    5'b00000: begin
                        WriteAddress<=7'd0;
                        ReadAddress<=7'd0;
                    end
                    
                    5'b00001: begin
                        WriteAddress<=7'd4;
                        ReadAddress<=7'd4;
                    end
                    
                    5'b00010: begin
                        WriteAddress<=7'd8;
                        ReadAddress<=7'd8;
                    end
                    
                    5'b00011: begin
                        WriteAddress<=7'd12;
                        ReadAddress<=7'd12;
                    end
                    
                    5'b00100: begin
                        WriteAddress<=7'd16;
                        ReadAddress<=7'd16;
                    end
                    
                    5'b00101: begin
                        WriteAddress<=7'd20;
                        ReadAddress<=7'd20;
                    end
                    
                    5'b00110: begin
                        WriteAddress<=7'd24;
                        ReadAddress<=7'd24;
                    end
                    
                    5'b00111: begin
                        WriteAddress<=7'd28;
                        ReadAddress<=7'd28;
                    end
                    
                    5'b01000: begin
                        WriteAddress<=7'd32;
                        ReadAddress<=7'd32;
                    end
                    
                    5'b01001: begin
                        WriteAddress<=7'd36;
                        ReadAddress<=7'd36;
                    end
                    
                    5'b01010: begin
                        WriteAddress<=7'd40;
                        ReadAddress<=7'd40;
                    end
                    
                    5'b01011: begin
                        WriteAddress<=7'd44;
                        ReadAddress<=7'd44;
                    end
                    
                    5'b01100: begin
                        WriteAddress<=7'd48;
                        ReadAddress<=7'd48;
                    end
                    
                    5'b01101: begin
                        WriteAddress<=7'd52;
                        ReadAddress<=7'd48;
                    end
                    
                    5'b01110: begin
                        WriteAddress<=7'd56;
                        ReadAddress<=7'd56;
                    end
                    
                    5'b01111: begin
                        WriteAddress<=7'd60;
                        ReadAddress<=7'd60;
                    end
                    
                    5'b10000: begin
                        WriteAddress<=7'd64;
                        ReadAddress<=7'd64;
                    end
                    
                    5'b10001: begin
                        WriteAddress<=7'd68;
                        ReadAddress<=7'd68;
                    end
                    
                    5'b10010: begin
                        WriteAddress<=7'd72;
                        ReadAddress<=7'd72;
                    end
                    
                    5'b10011: begin
                        WriteAddress<=7'd76;
                        ReadAddress<=7'd76;
                    end
                    
                    5'b10100: begin
                        WriteAddress<=7'd80;
                        ReadAddress<=7'd80;
                    end
                    
                    5'b10101: begin
                        WriteAddress<=7'd84;
                        ReadAddress<=7'd84;
                    end
                    
                    5'b10110: begin
                        WriteAddress<=7'd88;
                        ReadAddress<=7'd88;
                    end
                    
                    5'b10111: begin
                        WriteAddress<=7'd92;
                        ReadAddress<=7'd92;
                    end
                    
                    5'b11000: begin
                        WriteAddress<=7'd96;
                        ReadAddress<=7'd96;
                    end
                    
                    5'b11001: begin
                        WriteAddress<=7'd100;
                        ReadAddress<=7'd100;
                    end
                    
                    5'b11010: begin
                        WriteAddress<=7'd104;
                        ReadAddress<=7'd104;
                    end
                    
                    5'b11011: begin
                        WriteAddress<=7'd108;
                        ReadAddress<=7'd108;
                    end
                    
                    5'b11100: begin
                        WriteAddress<=7'd112;
                        ReadAddress<=7'd112;
                    end
                    
                    5'b11101: begin
                        WriteAddress<=7'd116;
                        ReadAddress<=7'd116;
                    end
                    
                    5'b11110: begin
                        WriteAddress<=7'd120;
                        ReadAddress<=7'd120;
                    end
                    
                    5'b11111: begin
                        WriteAddress<=7'd124;
                        ReadAddress<=7'd124;
                    end
                    
                    default: begin
                        WriteAddress<=7'd0;
                        ReadAddress<=7'd0;
                    end
                endcase
                end
            end
        else if(state==4'b0001)//write address and data keep for 2 cycle
            begin
                state<=4'b0010;
            end
        else if(state==4'b0010)
            begin
                write_en<=1'b0;
                read_en<=1'b1;
                rwControl<=1'b0;
                WriteAddress<=7'b0;
                state<=4'b0000;
                stop_reg<=1;
            end
end

endmodule
    
module compute_aux_write_aux2(
    input clk,
    input rst,
    input [254:0] data_in,
    input start,
    input [4:0] round,
    
    output  stop,
    output  [511:0] out
    //output [4:0] state_out
);

reg [6:0] WriteAddress, ReadAddress;
reg rwControl, read_en, write_en;
reg [511:0] data;
reg [3:0] state;
reg stop_reg;
wire [511:0] data_out;

assign out=data_out;
//assign state_out=state;
assign stop=stop_reg;


aux_bits aux 
(
  .clka(clk),    // input wire clka
  .ena(write_en),      // input wire ena
  .wea(rwControl),      // input wire [0 : 0] wea
  .addra(WriteAddress),  // input wire [6 : 0] addra
  .dina(data),    // input wire [511 : 0] dina
  .clkb(clk),    // input wire clkb
  .enb(read_en),      // input wire enb
  .addrb(ReadAddress),  // input wire [6 : 0] addrb
  .doutb(data_out)  // output wire [511 : 0] doutb
);
    
    
always@(posedge clk or negedge rst)
begin
    if(!rst)
        begin
            data<=512'b0;
            write_en<=1'b0;
            read_en<=1'b0;
            rwControl<=1'b0;
            state<=4'b0000;
            ReadAddress<=7'b0;
            WriteAddress<=7'b0;
        end
    else
        if(state==4'b0000)
            begin
                stop_reg<=0;
                if(start)
                begin

                    data<=512'b0;
                    state<=4'b0001;
                    rwControl<=1'b0;
                    write_en<=1'b0;
                    read_en<=1'b1;

                case(round)
                    5'b00000: begin
                        WriteAddress<=7'd0;
                        ReadAddress<=7'd0;
                    end
                    
                    5'b00001: begin
                        WriteAddress<=7'd4;
                        ReadAddress<=7'd4;
                    end
                    
                    5'b00010: begin
                        WriteAddress<=7'd8;
                        ReadAddress<=7'd8;
                    end
                    
                    5'b00011: begin
                        WriteAddress<=7'd12;
                        ReadAddress<=7'd12;
                    end
                    
                    5'b00100: begin
                        WriteAddress<=7'd16;
                        ReadAddress<=7'd16;
                    end
                    
                    5'b00101: begin
                        WriteAddress<=7'd20;
                        ReadAddress<=7'd20;
                    end
                    
                    5'b00110: begin
                        WriteAddress<=7'd24;
                        ReadAddress<=7'd24;
                    end
                    
                    5'b00111: begin
                        WriteAddress<=7'd28;
                        ReadAddress<=7'd28;
                    end
                    
                    5'b01000: begin
                        WriteAddress<=7'd32;
                        ReadAddress<=7'd32;
                    end
                    
                    5'b01001: begin
                        WriteAddress<=7'd36;
                        ReadAddress<=7'd36;
                    end
                    
                    5'b01010: begin
                        WriteAddress<=7'd40;
                        ReadAddress<=7'd40;
                    end
                    
                    5'b01011: begin
                        WriteAddress<=7'd44;
                        ReadAddress<=7'd44;
                    end
                    
                    5'b01100: begin
                        WriteAddress<=7'd48;
                        ReadAddress<=7'd48;
                    end
                    
                    5'b01101: begin
                        WriteAddress<=7'd52;
                        ReadAddress<=7'd48;
                    end
                    
                    5'b01110: begin
                        WriteAddress<=7'd56;
                        ReadAddress<=7'd56;
                    end
                    
                    5'b01111: begin
                        WriteAddress<=7'd60;
                        ReadAddress<=7'd60;
                    end
                    
                    5'b10000: begin
                        WriteAddress<=7'd64;
                        ReadAddress<=7'd64;
                    end
                    
                    5'b10001: begin
                        WriteAddress<=7'd68;
                        ReadAddress<=7'd68;
                    end
                    
                    5'b10010: begin
                        WriteAddress<=7'd72;
                        ReadAddress<=7'd72;
                    end
                    
                    5'b10011: begin
                        WriteAddress<=7'd76;
                        ReadAddress<=7'd76;
                    end
                    
                    5'b10100: begin
                        WriteAddress<=7'd80;
                        ReadAddress<=7'd80;
                    end
                    
                    5'b10101: begin
                        WriteAddress<=7'd84;
                        ReadAddress<=7'd84;
                    end
                    
                    5'b10110: begin
                        WriteAddress<=7'd88;
                        ReadAddress<=7'd88;
                    end
                    
                    5'b10111: begin
                        WriteAddress<=7'd92;
                        ReadAddress<=7'd92;
                    end
                    
                    5'b11000: begin
                        WriteAddress<=7'd96;
                        ReadAddress<=7'd96;
                    end
                    
                    5'b11001: begin
                        WriteAddress<=7'd100;
                        ReadAddress<=7'd100;
                    end
                    
                    5'b11010: begin
                        WriteAddress<=7'd104;
                        ReadAddress<=7'd104;
                    end
                    
                    5'b11011: begin
                        WriteAddress<=7'd108;
                        ReadAddress<=7'd108;
                    end
                    
                    5'b11100: begin
                        WriteAddress<=7'd112;
                        ReadAddress<=7'd112;
                    end
                    
                    5'b11101: begin
                        WriteAddress<=7'd116;
                        ReadAddress<=7'd116;
                    end
                    
                    5'b11110: begin
                        WriteAddress<=7'd120;
                        ReadAddress<=7'd120;
                    end
                    
                    5'b11111: begin
                        WriteAddress<=7'd124;
                        ReadAddress<=7'd124;
                    end
                    
                    default: begin
                        WriteAddress<=7'd0;
                        ReadAddress<=7'd0;
                    end
                endcase
                end
            end
        else if(state==4'b0001)//write address and data keep for 2 cycle
            begin
                data<={data_in, 1'b0, data_out[255:0]};
                read_en<=1'b0;
                write_en<=1'b1;
                rwControl<=1'b1;
                state<=4'b0010;
            end
        else if(state==4'b0010)
            begin
                write_en<=1'b0;
                read_en<=1'b1;
                rwControl<=1'b0;
                WriteAddress<=7'b0;
                state<=4'b0000;
                stop_reg<=1;
            end
end

endmodule    

module compute_aux_sm4_round(
    input clk,
    input rst,
    input [31:0] round_key_input1,
    input [31:0] round_key_input2,
    input start,
    
    output stop,
    output [3:0] state_out,
    output [254:0] test_out1,
    output [254:0] test_out2,
    output [511:0] inside_out1,
    output [511:0] inside_out2
    );
    wire [1019:0] aux_bits1, aux_bits2;
    reg [5:0] round;
    reg start1, start2, start3, start4;
    reg start5, start6, start7, start8;
    reg start9, start10;
    wire stop1, stop2, stop3, stop4;
    wire stop5, stop6, stop7, stop8;
    wire stop9, stop10;
    wire [254:0] xor_result1, xor_result2, xor_result3, xor_result4;
    wire [254:0] xor_result5, xor_result6, xor_result7, xor_result8;
    wire [511:0] inside_data1, inside_data2;
    reg [3:0] state;
    reg stop_reg;
    reg [254:0] final_xor_result1, final_xor_result2;
    reg dec;
    
    assign stop=stop_reg;
    assign state_out=state;
    assign test_out1=final_xor_result1;
    assign test_out2=final_xor_result2;
    assign inside_out1=inside_data1;
    assign inside_out2=inside_data2;
    
    compute_aux_bits CAB1(round_key_input1, aux_bits1);
    compute_aux_bits CAB2(round_key_input2, aux_bits2);
    
    compute_aux_read_tapes CART1(clk, rst, round, 2'b00, start1, 1'b0, xor_result1, stop1);
    compute_aux_read_tapes CART2(clk, rst, round, 2'b01, start2, 1'b0, xor_result2, stop2);
    compute_aux_read_tapes CART3(clk, rst, round, 2'b10, start3, 1'b0, xor_result3, stop3);
    compute_aux_read_tapes CART4(clk, rst, round, 2'b11, start4, 1'b0, xor_result4, stop4);
    
    compute_aux_write_aux1 CAWA1(clk, rst, final_xor_result1, start9, round, stop9, inside_data1);
    
    compute_aux_read_tapes CART5(clk, rst, round, 2'b00, start5, 1'b1, xor_result5, stop5);
    compute_aux_read_tapes CART6(clk, rst, round, 2'b01, start6, 1'b1, xor_result6, stop6);
    compute_aux_read_tapes CART7(clk, rst, round, 2'b10, start7, 1'b1, xor_result7, stop7);
    compute_aux_read_tapes CART8(clk, rst, round, 2'b11, start8, 1'b1, xor_result8, stop8);
    
    compute_aux_write_aux2 CAWA2(clk, rst, final_xor_result2, start10, round, stop10, inside_data2);
    always@(posedge clk or negedge rst)
    begin
        if(!rst)
            begin
                state<=4'b0000;
                stop_reg<=1'b0;
                final_xor_result1<=255'b0;
                final_xor_result2<=255'b0;
            end
        else
            begin
                if(state==4'b0000)
                    begin
                        stop_reg<=1'b0;
                        if(start)
                            begin
                                round<=5'b00000;
                                start1<=1'b0;
                                start2<=1'b0;
                                start3<=1'b0;
                                start4<=1'b0;
                                start5<=1'b0;
                                start6<=1'b0;
                                start7<=1'b0;
                                start8<=1'b0;
                                start9<=1'b0;
                                start9<=1'b0;
                                start10<=1'b0;
                                state<=4'b0001;
                                final_xor_result1<=255'b0;
                                final_xor_result2<=255'b0;
                                dec<=1'b0;
                            end
                    end
                else if(state==4'b0001)
                    begin
                        start1<=1'b1;
                        if(stop1)
                            begin
                                final_xor_result1<=final_xor_result1^xor_result1;
                                state<=4'b0010;
                                start1<=1'b0;
                            end
                    end
                    
                else if(state==4'b0010)
                    begin
                        start2<=1'b1;
                        if(stop2)
                            begin
                                final_xor_result1<=final_xor_result1^xor_result2;
                                state<=4'b0011;
                                start2<=1'b0;
                            end
                    end
                    
                else if(state==4'b0011)
                    begin
                        start3<=1'b1;
                        if(stop3)
                            begin
                                final_xor_result1<=final_xor_result1^xor_result3;
                                state<=4'b0100;
                                start3<=1'b0;
                            end
                    end
                    
                else if(state==4'b0100)
                    begin
                        start4<=1'b1;
                        if(stop4)
                            begin
                                final_xor_result1<=final_xor_result1^xor_result4;
                                state<=4'b0101;
                                start4<=1'b0;
                            end
                    end
                    
                else if(state==4'b0101)
                    begin
                        start9<=1'b1;
                        if(stop9)
                            begin
                                final_xor_result1<=255'b0;
                                state<=4'b0110;
                                start9<=1'b0;
                            end
                    end
                else if(state==4'b0110)
                    begin
                        start5<=1'b1;
                        if(stop5)
                            begin
                                final_xor_result2<=final_xor_result2^xor_result5;
                                state<=4'b0111;
                                start5<=1'b0;
                            end
                    end
                else if(state==4'b0111)
                    begin
                        start6<=1'b1;
                        if(stop6)
                            begin
                                final_xor_result2<=final_xor_result2^xor_result6;
                                state<=4'b1000;
                                start6<=1'b0;
                            end
                    end
                    
                else if(state==4'b1000)
                    begin
                        start7<=1'b1;
                        if(stop7)
                            begin
                                final_xor_result2<=final_xor_result2^xor_result7;
                                state<=4'b1001;
                                start7<=1'b0;
                            end
                    end
                    
                else if(state==4'b1001)
                    begin
                        start8<=1'b1;
                        if(stop8)
                            begin
                                final_xor_result2<=final_xor_result2^xor_result8;
                                state<=4'b1010;
                                start8<=1'b0;
                            end
                    end
                else if(state==4'b1010)
                    begin
                        start10<=1'b1;
                        if(stop10)
                            begin
                                final_xor_result2<=255'b0;
                                state<=4'b0000;
                                stop_reg<=1'b1;
                                start10<=1'b0;
                            end
                        
                    end
            end
    end
    
endmodule

module Get_Read_Address(
    input [4:0] round,
    input [1:0] k,
    output  reg [10:0] ReadAddress
);
    always@(*)
    begin
                    case(round)
                        5'b00000: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd0;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd1;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd2;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd3;
                                end
                            endcase
                        end
                        
                        5'b00001: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd4;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd5;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd6;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd7;
                                end
                            endcase
                        end
                        
                        5'b00010: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd8;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd9;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd10;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd11;
                                end
                            endcase
                        end
                        
                        5'b00011: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd12;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd13;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd14;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd15;
                                end
                            endcase
                        end
                        
                        5'b00100: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd16;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd17;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd18;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd19;
                                end
                            endcase
                        end
                        
                        5'b00101: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd20;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd21;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd22;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd23;
                                end
                            endcase
                        end
                        
                        5'b00110: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd24;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd25;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd26;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd27;
                                end
                            endcase
                        end
                        
                        5'b00111: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd28;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd29;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd30;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd31;
                                end
                            endcase
                        end
                        
                        5'b01000: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd32;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd33;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd34;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd35;
                                end
                            endcase
                        end
                        
                        5'b01001: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd36;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd37;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd38;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd39;
                                end
                            endcase
                        end
                        
                        5'b01010: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd40;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd41;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd42;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd43;
                                end
                            endcase
                        end
                        
                        5'b01011: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd44;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd45;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd46;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd47;
                                end
                            endcase
                        end
                        
                        5'b01100: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd48;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd49;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd50;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd51;
                                end
                            endcase
                        end
                        
                        5'b01101: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd52;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd53;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd54;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd55;
                                end
                            endcase
                        end
                        
                        5'b01110: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd56;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd57;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd58;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd59;
                                end
                            endcase
                        end
                        
                        5'b01111: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd60;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd61;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd62;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd63;
                                end
                            endcase
                        end
                        
                        5'b10000: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd64;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd65;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd66;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd67;
                                end
                            endcase
                        end
                        
                        5'b10001: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd68;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd69;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd70;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd71;
                                end
                            endcase
                        end
                        
                        5'b10010: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd72;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd73;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd74;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd75;
                                end
                            endcase
                        end
                        
                        5'b10011: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd76;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd77;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd78;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd79;
                                end
                            endcase
                        end
                        
                        5'b10100: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd80;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd81;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd82;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd83;
                                end
                            endcase
                        end
                        
                        5'b10101: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd84;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd85;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd86;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd87;
                                end
                            endcase
                        end
                        
                        5'b10110: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd88;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd89;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd90;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd91;
                                end
                            endcase
                        end
                        
                        5'b10111: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd92;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd93;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd94;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd95;
                                end
                            endcase
                        end
                        
                        5'b11000: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd96;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd97;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd98;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd99;
                                end
                            endcase
                        end
                        
                        5'b11001: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd100;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd101;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd102;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd103;
                                end
                            endcase
                        end
                        
                        5'b11010: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd104;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd105;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd106;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd107;
                                end
                            endcase
                        end
                        
                        5'b11011: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd108;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd109;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd110;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd111;
                                end
                            endcase
                        end
                        
                        5'b11100: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd112;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd113;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd114;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd115;
                                end
                            endcase
                        end
                        
                        5'b11101: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd116;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd117;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd118;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd119;
                                end
                            endcase
                        end
                        
                        5'b11110: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd120;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd121;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd122;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd123;
                                end
                            endcase
                        end
                        
                        5'b11111: begin
                            case(k)
                                2'b00: begin
                                    ReadAddress<=11'd124;
                                end
                                
                                2'b01: begin
                                    ReadAddress<=11'd125;
                                end
                                
                                2'b10: begin
                                    ReadAddress<=11'd126;
                                end
                                
                                2'b11: begin
                                    ReadAddress<=11'd127;
                                end
                            endcase
                        end
                        
                        
                        default: begin
                            ReadAddress<=11'b0;
                        end
                    endcase
                end
endmodule

module Get_Write_Address(
    input [4:0] round,
    output reg [6:0] WriteAddress
);
    always@(*)
    begin
        case(round)
                    5'b00000: begin
                        WriteAddress<=7'd0;

                    end
                    
                    5'b00001: begin
                        WriteAddress<=7'd4;

                    end
                    
                    5'b00010: begin
                        WriteAddress<=7'd8;

                    end
                    
                    5'b00011: begin
                        WriteAddress<=7'd12;

                    end
                    
                    5'b00100: begin
                        WriteAddress<=7'd16;

                    end
                    
                    5'b00101: begin
                        WriteAddress<=7'd20;

                    end
                    
                    5'b00110: begin
                        WriteAddress<=7'd24;

                    end
                    
                    5'b00111: begin
                        WriteAddress<=7'd28;

                    end
                    
                    5'b01000: begin
                        WriteAddress<=7'd32;

                    end
                    
                    5'b01001: begin
                        WriteAddress<=7'd36;

                    end
                    
                    5'b01010: begin
                        WriteAddress<=7'd40;

                    end
                    
                    5'b01011: begin
                        WriteAddress<=7'd44;

                    end
                    
                    5'b01100: begin
                        WriteAddress<=7'd48;

                    end
                    
                    5'b01101: begin
                        WriteAddress<=7'd52;

                    end
                    
                    5'b01110: begin
                        WriteAddress<=7'd56;

                    end
                    
                    5'b01111: begin
                        WriteAddress<=7'd60;

                    end
                    
                    5'b10000: begin
                        WriteAddress<=7'd64;

                    end
                    
                    5'b10001: begin
                        WriteAddress<=7'd68;

                    end
                    
                    5'b10010: begin
                        WriteAddress<=7'd72;

                    end
                    
                    5'b10011: begin
                        WriteAddress<=7'd76;

                    end
                    
                    5'b10100: begin
                        WriteAddress<=7'd80;

                    end
                    
                    5'b10101: begin
                        WriteAddress<=7'd84;

                    end
                    
                    5'b10110: begin
                        WriteAddress<=7'd88;

                    end
                    
                    5'b10111: begin
                        WriteAddress<=7'd92;

                    end
                    
                    5'b11000: begin
                        WriteAddress<=7'd96;

                    end
                    
                    5'b11001: begin
                        WriteAddress<=7'd100;

                    end
                    
                    5'b11010: begin
                        WriteAddress<=7'd104;

                    end
                    
                    5'b11011: begin
                        WriteAddress<=7'd108;

                    end
                    
                    5'b11100: begin
                        WriteAddress<=7'd112;

                    end
                    
                    5'b11101: begin
                        WriteAddress<=7'd116;

                    end
                    
                    5'b11110: begin
                        WriteAddress<=7'd120;

                    end
                    
                    5'b11111: begin
                        WriteAddress<=7'd124;

                    end
                    
                    default: begin
                        WriteAddress<=7'd0;

                    end
                endcase
    end
endmodule


module Get_RoundKey_xor(
    input [4:0] round,
    input [1:0] t,
    
    output reg [31:0] xor_result
);

    always@(*)
    begin
        case(round)
                    5'b00000: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h3de5e1fc;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h7b2b5dc1;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h92b2aa38;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h643224e;
                            end
                            
                        endcase
                    end
                    
                    5'b00001: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h6c56f7eb;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h2fab1496;
                            end
                            
                            2'b10: begin
                                xor_result<=32'ha41cf8c4;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h8181d279;
                            end
                            
                        endcase
                    end
                    
                    5'b00010: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h2057026a;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h1176a667;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hcd47b36c;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hddf25360;
                            end
                            
                        endcase
                    end
                    
                    5'b00011: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h1c5deb0;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hef4d89ab;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h45fd05b;
                            end
                            
                            2'b11: begin
                                xor_result<=32'ha89b424b;
                            end
                            
                        endcase
                    end
                    
                    5'b00100: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h16bcd21b;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hce1ebaee;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h4e0a3511;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h3415c9a4;
                            end
                            
                        endcase
                    end
                    
                    5'b00101: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hc1a46603;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hbce01f23;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h1ea316cf;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hccd7b405;
                            end
                            
                        endcase
                    end
                    
                    5'b00110: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'ha73fa2f3;
                            end
                            
                            2'b01: begin
                                xor_result<=32'he5345a19;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h7960d0ca;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h45ee96aa;
                            end
                            
                        endcase
                    end
                    
                    5'b00111: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hf01d33bb;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h49d74b4c;
                            end
                            
                            2'b10: begin
                                xor_result<=32'ha3b0eafd;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h507fab7c;
                            end
                            
                        endcase
                    end
                    
                    5'b01000: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hbf1379dd;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h84de7bbb;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h2866e5cf;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hd7aa51be;
                            end
                            
                        endcase
                    end
                    
                    5'b01001: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h91401c1f;
                            end
                            
                            2'b01: begin
                                xor_result<=32'he8d24309;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h3355ce0a;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h231b0a58;
                            end
                            
                        endcase
                    end
                    
                    5'b01010: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hd59a1b06;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hf250c90e;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h217bc79a;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hfaeba03e;
                            end
                            
                        endcase
                    end
                    
                    5'b01011: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h5f6e46fd;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h27e9596;
                            end
                            
                            2'b10: begin
                                xor_result<=32'heba31b1c;
                            end
                            
                            2'b11: begin
                                xor_result<=32'heec08c37;
                            end
                            
                        endcase
                    end
                    
                    5'b01100: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h75748331;
                            end
                            
                            2'b01: begin    
                                xor_result<=32'hc19cbf2a;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hc3a33046;
                            end
                            
                            2'b11: begin
                                xor_result<=32'ha92dd47b;
                            end
                            
                        endcase
                    end
                    
                    5'b01101: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h7d22bbdb;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h574ab713;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hbb8c307d;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h39fc6ab9;
                            end
                            
                        endcase
                    end
                    
                    5'b01110: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hde5d3c13;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h119a55b2;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hecf44a3a;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hfb4a8508;
                            end
                            
                        endcase
                    end
                    
                    5'b01111: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hf4663106;
                            end 
                            
                            2'b01: begin
                                xor_result<=32'ha15d2e81;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h7d3c7838;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h74cdc970;
                            end
                            
                        endcase
                    end
                    
                    5'b10000: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h195470c6;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hcff48241;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h4521807a;
                            end
                            
                            2'b11: begin
                                xor_result<=32'headfbf4c;
                            end
                            
                        endcase
                    end
                    
                    5'b10001: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h57576fd5;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hcfdd6a44;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h426dd39c;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hb5773126;
                            end
                            
                        endcase
                    end
                    
                    5'b10010: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hc4c14f7d;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h500931f8;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hd3631beb;
                            end
                            
                            2'b11: begin
                                xor_result<=32'ha7d13369;
                            end
                            
                        endcase
                    end
                    
                    5'b10011: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hafa50ae3;
                            end
                            
                            2'b01: begin
                                xor_result<=32'he790bce2;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h17cc667;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h7d98c09e;
                            end
                            
                        endcase
                    end
                    
                    5'b10100: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h262a346;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h58aaa666;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hc3e7fc7a;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h195df60f;
                            end
                            
                        endcase
                    end
                    
                    5'b10101: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hae4c3a95;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h6f30667b;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h79fe6353;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hab03232c;
                            end
                            
                        endcase
                    end
                    
                    5'b10110: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h86f86092;
                            end 
                            
                            2'b01: begin
                                xor_result<=32'h383a261b;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hb4a92ab8;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h31994ef8;
                            end
                            
                        endcase
                    end
                    
                    5'b10111: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hca77943;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hd9031460;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hb1abd299;
                            end
                            
                            2'b11: begin
                                xor_result<=32'ha2274721;
                            end
                            
                        endcase
                    end
                    
                    5'b11000: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h74fa9a68;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h6209b14;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hd6e66bf9;
                            end
                            
                            2'b11: begin
                                xor_result<=32'ha0666b88;
                            end
                            
                        endcase
                    end
                    
                    5'b11001: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hb40756d2;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h808b80b;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h707d95f3;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h2a64a90d;
                            end
                            
                        endcase
                    end
                    
                    5'b11010: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hfed3523a;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h49e00bcc;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hae2bdeb0;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h271d2214;
                            end
                            
                        endcase
                    end
                    
                    5'b11011: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h167c8ce7;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h6f7259cd;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h7b1bde1f;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h5bb4348d;
                            end
                            
                        endcase
                    end
                    
                    5'b11100: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h2a7435bd;
                            end
                            
                            2'b01: begin
                                xor_result<=32'he0ac131b;
                            end
                            
                            2'b10: begin
                                xor_result<=32'hdf03aa88;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h2161d1f3;
                            end
                            
                        endcase
                    end
                    
                    5'b11101: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hbe090b8e;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h86af96ad;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h9a6a362c;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h33f93779;
                            end
                            
                        endcase
                    end
                    
                    5'b11110: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'h82ff33f6;
                            end
                            
                            2'b01: begin
                                xor_result<=32'h4dbedabb;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h69414641;
                            end
                            
                            2'b11: begin
                                xor_result<=32'h3d82ab79;
                            end
                            
                        endcase
                    end
                    
                    5'b11111: begin
                        case (t)
                            2'b00: begin
                                xor_result<=32'hc7cd2987;
                            end
                            
                            2'b01: begin
                                xor_result<=32'hb13adfa0;
                            end
                            
                            2'b10: begin
                                xor_result<=32'h99fe91b5;
                            end
                            
                            2'b11: begin
                                xor_result<=32'hfbc69655;
                            end
                            
                        endcase
                    end
                    
                    default: begin
                        xor_result<=32'h0;
                    end
        endcase
    end
    
endmodule


module Get_Plaintext(
    input [5:0] index,
    output reg [31:0] plaintext
);

    
    always@(*)
    begin
        case(index)
            6'd0: begin
                plaintext<=32'h2f5b89a;
            end
            
            6'd1: begin
                plaintext<=32'haf493824;
            end
            
            6'd2: begin
                plaintext<=32'h71e9a340;
            end
            
            6'd3: begin
                plaintext<=32'h19bce013;
            end
            
            6'd4: begin
                plaintext<=32'h2794dec2;
            end
            
            6'd5: begin
                plaintext<=32'hde6a5985;
            end
            
            6'd6: begin
                plaintext<=32'hcf31974a;
            end
            
            6'd7: begin
                plaintext<=32'h56e9f864;
            end
            
            6'd8: begin
                plaintext<=32'h871cbf37;
            end
            
            6'd9: begin
                plaintext<=32'h758d14f8;
            end
            
            6'd10: begin
                plaintext<=32'hd372e9cc;
            end
            
            6'd11: begin
                plaintext<=32'hcddfbbaf;
            end
            
            6'd12: begin
                plaintext<=32'h6c32767a;
            end
            
            6'd13: begin
                plaintext<=32'h2aadb87b;
            end
            
            6'd14: begin
                plaintext<=32'ha8c16571;
            end
            
            6'd15: begin
                plaintext<=32'h71b39269;
            end
            
            6'd16: begin
                plaintext<=32'h39a2f357;
            end
            
            6'd17: begin
                plaintext<=32'h9c1ba044;
            end
            
            6'd18: begin
                plaintext<=32'hb13dd32c;
            end
            
            6'd19: begin
                plaintext<=32'h476d2161;
            end
            
            6'd20: begin
                plaintext<=32'hf6dfc65a;
            end
            
            6'd21: begin
                plaintext<=32'h48ccb222;
            end
            
            6'd22: begin
                plaintext<=32'hd4b15e06;
            end
            
            6'd23: begin
                plaintext<=32'h7b9373d0;
            end
            
            6'd24: begin
                plaintext<=32'h582ffd19;
            end
            
            6'd25: begin
                plaintext<=32'h3bd028ff;
            end
            
            6'd26: begin
                plaintext<=32'h9247e362;
            end
            
            6'd27: begin
                plaintext<=32'h82575bda;
            end
            
            6'd28: begin
                plaintext<=32'h78ebf11;
            end
            
            6'd29: begin
                plaintext<=32'h277507b7;
            end
            
            6'd30: begin
                plaintext<=32'h1aa0adf8;
            end
            
            6'd31: begin
                plaintext<=32'hcfd5bf01;
            end
            
            6'd32: begin
                plaintext<=32'h375bf876;
            end
            
            6'd33: begin
                plaintext<=32'h3a0eb9b2;
            end
            
            6'd34: begin
                plaintext<=32'h43bcecb4;
            end
            
            6'd35: begin
                plaintext<=32'hadc80985;
            end
            
            default: begin
                plaintext<=32'h2f5b89a;
            end
        endcase
    end
endmodule

