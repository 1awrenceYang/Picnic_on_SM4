module w_ram_from_sign
(
	input wire sys_clk,
	input wire sys_rst_n,
	input [19584-1:0] sigma_out,
    input wire w_ram_from_sign_start,
	output reg [7:0] data,
	output[14:0] address,
	output reg wea,
	output reg w_ram_from_sign_end
);

wire[14:0] full_number=2448;

wire[7:0] uart_rx_data;


reg[14:0] counter;

reg[2:0] state;

assign address = counter;

wire [7:0]sigma_out_list[2447:0];
assign {sigma_out_list[0],sigma_out_list[1],sigma_out_list[2],sigma_out_list[3],sigma_out_list[4],sigma_out_list[5],sigma_out_list[6],sigma_out_list[7],sigma_out_list[8],sigma_out_list[9],sigma_out_list[10],sigma_out_list[11],sigma_out_list[12],sigma_out_list[13],sigma_out_list[14],sigma_out_list[15],sigma_out_list[16],sigma_out_list[17],sigma_out_list[18],sigma_out_list[19],sigma_out_list[20],sigma_out_list[21],sigma_out_list[22],sigma_out_list[23],sigma_out_list[24],sigma_out_list[25],sigma_out_list[26],sigma_out_list[27],sigma_out_list[28],sigma_out_list[29],sigma_out_list[30],sigma_out_list[31],sigma_out_list[32],sigma_out_list[33],sigma_out_list[34],sigma_out_list[35],sigma_out_list[36],sigma_out_list[37],sigma_out_list[38],sigma_out_list[39],sigma_out_list[40],sigma_out_list[41],sigma_out_list[42],sigma_out_list[43],sigma_out_list[44],sigma_out_list[45],sigma_out_list[46],sigma_out_list[47],sigma_out_list[48],sigma_out_list[49],sigma_out_list[50],sigma_out_list[51],sigma_out_list[52],sigma_out_list[53],sigma_out_list[54],sigma_out_list[55],sigma_out_list[56],sigma_out_list[57],sigma_out_list[58],sigma_out_list[59],sigma_out_list[60],sigma_out_list[61],sigma_out_list[62],sigma_out_list[63],sigma_out_list[64],sigma_out_list[65],sigma_out_list[66],sigma_out_list[67],sigma_out_list[68],sigma_out_list[69],sigma_out_list[70],sigma_out_list[71],sigma_out_list[72],sigma_out_list[73],sigma_out_list[74],sigma_out_list[75],sigma_out_list[76],sigma_out_list[77],sigma_out_list[78],sigma_out_list[79],sigma_out_list[80],sigma_out_list[81],sigma_out_list[82],sigma_out_list[83],sigma_out_list[84],sigma_out_list[85],sigma_out_list[86],sigma_out_list[87],sigma_out_list[88],sigma_out_list[89],sigma_out_list[90],sigma_out_list[91],sigma_out_list[92],sigma_out_list[93],sigma_out_list[94],sigma_out_list[95],sigma_out_list[96],sigma_out_list[97],sigma_out_list[98],sigma_out_list[99],sigma_out_list[100],sigma_out_list[101],sigma_out_list[102],sigma_out_list[103],sigma_out_list[104],sigma_out_list[105],sigma_out_list[106],sigma_out_list[107],sigma_out_list[108],sigma_out_list[109],sigma_out_list[110],sigma_out_list[111],sigma_out_list[112],sigma_out_list[113],sigma_out_list[114],sigma_out_list[115],sigma_out_list[116],sigma_out_list[117],sigma_out_list[118],sigma_out_list[119],sigma_out_list[120],sigma_out_list[121],sigma_out_list[122],sigma_out_list[123],sigma_out_list[124],sigma_out_list[125],sigma_out_list[126],sigma_out_list[127],sigma_out_list[128],sigma_out_list[129],sigma_out_list[130],sigma_out_list[131],sigma_out_list[132],sigma_out_list[133],sigma_out_list[134],sigma_out_list[135],sigma_out_list[136],sigma_out_list[137],sigma_out_list[138],sigma_out_list[139],sigma_out_list[140],sigma_out_list[141],sigma_out_list[142],sigma_out_list[143],sigma_out_list[144],sigma_out_list[145],sigma_out_list[146],sigma_out_list[147],sigma_out_list[148],sigma_out_list[149],sigma_out_list[150],sigma_out_list[151],sigma_out_list[152],sigma_out_list[153],sigma_out_list[154],sigma_out_list[155],sigma_out_list[156],sigma_out_list[157],sigma_out_list[158],sigma_out_list[159],sigma_out_list[160],sigma_out_list[161],sigma_out_list[162],sigma_out_list[163],sigma_out_list[164],sigma_out_list[165],sigma_out_list[166],sigma_out_list[167],sigma_out_list[168],sigma_out_list[169],sigma_out_list[170],sigma_out_list[171],sigma_out_list[172],sigma_out_list[173],sigma_out_list[174],sigma_out_list[175],sigma_out_list[176],sigma_out_list[177],sigma_out_list[178],sigma_out_list[179],sigma_out_list[180],sigma_out_list[181],sigma_out_list[182],sigma_out_list[183],sigma_out_list[184],sigma_out_list[185],sigma_out_list[186],sigma_out_list[187],sigma_out_list[188],sigma_out_list[189],sigma_out_list[190],sigma_out_list[191],sigma_out_list[192],sigma_out_list[193],sigma_out_list[194],sigma_out_list[195],sigma_out_list[196],sigma_out_list[197],sigma_out_list[198],sigma_out_list[199],sigma_out_list[200],sigma_out_list[201],sigma_out_list[202],sigma_out_list[203],sigma_out_list[204],sigma_out_list[205],sigma_out_list[206],sigma_out_list[207],sigma_out_list[208],sigma_out_list[209],sigma_out_list[210],sigma_out_list[211],sigma_out_list[212],sigma_out_list[213],sigma_out_list[214],sigma_out_list[215],sigma_out_list[216],sigma_out_list[217],sigma_out_list[218],sigma_out_list[219],sigma_out_list[220],sigma_out_list[221],sigma_out_list[222],sigma_out_list[223],sigma_out_list[224],sigma_out_list[225],sigma_out_list[226],sigma_out_list[227],sigma_out_list[228],sigma_out_list[229],sigma_out_list[230],sigma_out_list[231],sigma_out_list[232],sigma_out_list[233],sigma_out_list[234],sigma_out_list[235],sigma_out_list[236],sigma_out_list[237],sigma_out_list[238],sigma_out_list[239],sigma_out_list[240],sigma_out_list[241],sigma_out_list[242],sigma_out_list[243],sigma_out_list[244],sigma_out_list[245],sigma_out_list[246],sigma_out_list[247],sigma_out_list[248],sigma_out_list[249],sigma_out_list[250],sigma_out_list[251],sigma_out_list[252],sigma_out_list[253],sigma_out_list[254],sigma_out_list[255],sigma_out_list[256],sigma_out_list[257],sigma_out_list[258],sigma_out_list[259],sigma_out_list[260],sigma_out_list[261],sigma_out_list[262],sigma_out_list[263],sigma_out_list[264],sigma_out_list[265],sigma_out_list[266],sigma_out_list[267],sigma_out_list[268],sigma_out_list[269],sigma_out_list[270],sigma_out_list[271],sigma_out_list[272],sigma_out_list[273],sigma_out_list[274],sigma_out_list[275],sigma_out_list[276],sigma_out_list[277],sigma_out_list[278],sigma_out_list[279],sigma_out_list[280],sigma_out_list[281],sigma_out_list[282],sigma_out_list[283],sigma_out_list[284],sigma_out_list[285],sigma_out_list[286],sigma_out_list[287],sigma_out_list[288],sigma_out_list[289],sigma_out_list[290],sigma_out_list[291],sigma_out_list[292],sigma_out_list[293],sigma_out_list[294],sigma_out_list[295],sigma_out_list[296],sigma_out_list[297],sigma_out_list[298],sigma_out_list[299],sigma_out_list[300],sigma_out_list[301],sigma_out_list[302],sigma_out_list[303],sigma_out_list[304],sigma_out_list[305],sigma_out_list[306],sigma_out_list[307],sigma_out_list[308],sigma_out_list[309],sigma_out_list[310],sigma_out_list[311],sigma_out_list[312],sigma_out_list[313],sigma_out_list[314],sigma_out_list[315],sigma_out_list[316],sigma_out_list[317],sigma_out_list[318],sigma_out_list[319],sigma_out_list[320],sigma_out_list[321],sigma_out_list[322],sigma_out_list[323],sigma_out_list[324],sigma_out_list[325],sigma_out_list[326],sigma_out_list[327],sigma_out_list[328],sigma_out_list[329],sigma_out_list[330],sigma_out_list[331],sigma_out_list[332],sigma_out_list[333],sigma_out_list[334],sigma_out_list[335],sigma_out_list[336],sigma_out_list[337],sigma_out_list[338],sigma_out_list[339],sigma_out_list[340],sigma_out_list[341],sigma_out_list[342],sigma_out_list[343],sigma_out_list[344],sigma_out_list[345],sigma_out_list[346],sigma_out_list[347],sigma_out_list[348],sigma_out_list[349],sigma_out_list[350],sigma_out_list[351],sigma_out_list[352],sigma_out_list[353],sigma_out_list[354],sigma_out_list[355],sigma_out_list[356],sigma_out_list[357],sigma_out_list[358],sigma_out_list[359],sigma_out_list[360],sigma_out_list[361],sigma_out_list[362],sigma_out_list[363],sigma_out_list[364],sigma_out_list[365],sigma_out_list[366],sigma_out_list[367],sigma_out_list[368],sigma_out_list[369],sigma_out_list[370],sigma_out_list[371],sigma_out_list[372],sigma_out_list[373],sigma_out_list[374],sigma_out_list[375],sigma_out_list[376],sigma_out_list[377],sigma_out_list[378],sigma_out_list[379],sigma_out_list[380],sigma_out_list[381],sigma_out_list[382],sigma_out_list[383],sigma_out_list[384],sigma_out_list[385],sigma_out_list[386],sigma_out_list[387],sigma_out_list[388],sigma_out_list[389],sigma_out_list[390],sigma_out_list[391],sigma_out_list[392],sigma_out_list[393],sigma_out_list[394],sigma_out_list[395],sigma_out_list[396],sigma_out_list[397],sigma_out_list[398],sigma_out_list[399],sigma_out_list[400],sigma_out_list[401],sigma_out_list[402],sigma_out_list[403],sigma_out_list[404],sigma_out_list[405],sigma_out_list[406],sigma_out_list[407],sigma_out_list[408],sigma_out_list[409],sigma_out_list[410],sigma_out_list[411],sigma_out_list[412],sigma_out_list[413],sigma_out_list[414],sigma_out_list[415],sigma_out_list[416],sigma_out_list[417],sigma_out_list[418],sigma_out_list[419],sigma_out_list[420],sigma_out_list[421],sigma_out_list[422],sigma_out_list[423],sigma_out_list[424],sigma_out_list[425],sigma_out_list[426],sigma_out_list[427],sigma_out_list[428],sigma_out_list[429],sigma_out_list[430],sigma_out_list[431],sigma_out_list[432],sigma_out_list[433],sigma_out_list[434],sigma_out_list[435],sigma_out_list[436],sigma_out_list[437],sigma_out_list[438],sigma_out_list[439],sigma_out_list[440],sigma_out_list[441],sigma_out_list[442],sigma_out_list[443],sigma_out_list[444],sigma_out_list[445],sigma_out_list[446],sigma_out_list[447],sigma_out_list[448],sigma_out_list[449],sigma_out_list[450],sigma_out_list[451],sigma_out_list[452],sigma_out_list[453],sigma_out_list[454],sigma_out_list[455],sigma_out_list[456],sigma_out_list[457],sigma_out_list[458],sigma_out_list[459],sigma_out_list[460],sigma_out_list[461],sigma_out_list[462],sigma_out_list[463],sigma_out_list[464],sigma_out_list[465],sigma_out_list[466],sigma_out_list[467],sigma_out_list[468],sigma_out_list[469],sigma_out_list[470],sigma_out_list[471],sigma_out_list[472],sigma_out_list[473],sigma_out_list[474],sigma_out_list[475],sigma_out_list[476],sigma_out_list[477],sigma_out_list[478],sigma_out_list[479],sigma_out_list[480],sigma_out_list[481],sigma_out_list[482],sigma_out_list[483],sigma_out_list[484],sigma_out_list[485],sigma_out_list[486],sigma_out_list[487],sigma_out_list[488],sigma_out_list[489],sigma_out_list[490],sigma_out_list[491],sigma_out_list[492],sigma_out_list[493],sigma_out_list[494],sigma_out_list[495],sigma_out_list[496],sigma_out_list[497],sigma_out_list[498],sigma_out_list[499],sigma_out_list[500],sigma_out_list[501],sigma_out_list[502],sigma_out_list[503],sigma_out_list[504],sigma_out_list[505],sigma_out_list[506],sigma_out_list[507],sigma_out_list[508],sigma_out_list[509],sigma_out_list[510],sigma_out_list[511],sigma_out_list[512],sigma_out_list[513],sigma_out_list[514],sigma_out_list[515],sigma_out_list[516],sigma_out_list[517],sigma_out_list[518],sigma_out_list[519],sigma_out_list[520],sigma_out_list[521],sigma_out_list[522],sigma_out_list[523],sigma_out_list[524],sigma_out_list[525],sigma_out_list[526],sigma_out_list[527],sigma_out_list[528],sigma_out_list[529],sigma_out_list[530],sigma_out_list[531],sigma_out_list[532],sigma_out_list[533],sigma_out_list[534],sigma_out_list[535],sigma_out_list[536],sigma_out_list[537],sigma_out_list[538],sigma_out_list[539],sigma_out_list[540],sigma_out_list[541],sigma_out_list[542],sigma_out_list[543],sigma_out_list[544],sigma_out_list[545],sigma_out_list[546],sigma_out_list[547],sigma_out_list[548],sigma_out_list[549],sigma_out_list[550],sigma_out_list[551],sigma_out_list[552],sigma_out_list[553],sigma_out_list[554],sigma_out_list[555],sigma_out_list[556],sigma_out_list[557],sigma_out_list[558],sigma_out_list[559],sigma_out_list[560],sigma_out_list[561],sigma_out_list[562],sigma_out_list[563],sigma_out_list[564],sigma_out_list[565],sigma_out_list[566],sigma_out_list[567],sigma_out_list[568],sigma_out_list[569],sigma_out_list[570],sigma_out_list[571],sigma_out_list[572],sigma_out_list[573],sigma_out_list[574],sigma_out_list[575],sigma_out_list[576],sigma_out_list[577],sigma_out_list[578],sigma_out_list[579],sigma_out_list[580],sigma_out_list[581],sigma_out_list[582],sigma_out_list[583],sigma_out_list[584],sigma_out_list[585],sigma_out_list[586],sigma_out_list[587],sigma_out_list[588],sigma_out_list[589],sigma_out_list[590],sigma_out_list[591],sigma_out_list[592],sigma_out_list[593],sigma_out_list[594],sigma_out_list[595],sigma_out_list[596],sigma_out_list[597],sigma_out_list[598],sigma_out_list[599],sigma_out_list[600],sigma_out_list[601],sigma_out_list[602],sigma_out_list[603],sigma_out_list[604],sigma_out_list[605],sigma_out_list[606],sigma_out_list[607],sigma_out_list[608],sigma_out_list[609],sigma_out_list[610],sigma_out_list[611],sigma_out_list[612],sigma_out_list[613],sigma_out_list[614],sigma_out_list[615],sigma_out_list[616],sigma_out_list[617],sigma_out_list[618],sigma_out_list[619],sigma_out_list[620],sigma_out_list[621],sigma_out_list[622],sigma_out_list[623],sigma_out_list[624],sigma_out_list[625],sigma_out_list[626],sigma_out_list[627],sigma_out_list[628],sigma_out_list[629],sigma_out_list[630],sigma_out_list[631],sigma_out_list[632],sigma_out_list[633],sigma_out_list[634],sigma_out_list[635],sigma_out_list[636],sigma_out_list[637],sigma_out_list[638],sigma_out_list[639],sigma_out_list[640],sigma_out_list[641],sigma_out_list[642],sigma_out_list[643],sigma_out_list[644],sigma_out_list[645],sigma_out_list[646],sigma_out_list[647],sigma_out_list[648],sigma_out_list[649],sigma_out_list[650],sigma_out_list[651],sigma_out_list[652],sigma_out_list[653],sigma_out_list[654],sigma_out_list[655],sigma_out_list[656],sigma_out_list[657],sigma_out_list[658],sigma_out_list[659],sigma_out_list[660],sigma_out_list[661],sigma_out_list[662],sigma_out_list[663],sigma_out_list[664],sigma_out_list[665],sigma_out_list[666],sigma_out_list[667],sigma_out_list[668],sigma_out_list[669],sigma_out_list[670],sigma_out_list[671],sigma_out_list[672],sigma_out_list[673],sigma_out_list[674],sigma_out_list[675],sigma_out_list[676],sigma_out_list[677],sigma_out_list[678],sigma_out_list[679],sigma_out_list[680],sigma_out_list[681],sigma_out_list[682],sigma_out_list[683],sigma_out_list[684],sigma_out_list[685],sigma_out_list[686],sigma_out_list[687],sigma_out_list[688],sigma_out_list[689],sigma_out_list[690],sigma_out_list[691],sigma_out_list[692],sigma_out_list[693],sigma_out_list[694],sigma_out_list[695],sigma_out_list[696],sigma_out_list[697],sigma_out_list[698],sigma_out_list[699],sigma_out_list[700],sigma_out_list[701],sigma_out_list[702],sigma_out_list[703],sigma_out_list[704],sigma_out_list[705],sigma_out_list[706],sigma_out_list[707],sigma_out_list[708],sigma_out_list[709],sigma_out_list[710],sigma_out_list[711],sigma_out_list[712],sigma_out_list[713],sigma_out_list[714],sigma_out_list[715],sigma_out_list[716],sigma_out_list[717],sigma_out_list[718],sigma_out_list[719],sigma_out_list[720],sigma_out_list[721],sigma_out_list[722],sigma_out_list[723],sigma_out_list[724],sigma_out_list[725],sigma_out_list[726],sigma_out_list[727],sigma_out_list[728],sigma_out_list[729],sigma_out_list[730],sigma_out_list[731],sigma_out_list[732],sigma_out_list[733],sigma_out_list[734],sigma_out_list[735],sigma_out_list[736],sigma_out_list[737],sigma_out_list[738],sigma_out_list[739],sigma_out_list[740],sigma_out_list[741],sigma_out_list[742],sigma_out_list[743],sigma_out_list[744],sigma_out_list[745],sigma_out_list[746],sigma_out_list[747],sigma_out_list[748],sigma_out_list[749],sigma_out_list[750],sigma_out_list[751],sigma_out_list[752],sigma_out_list[753],sigma_out_list[754],sigma_out_list[755],sigma_out_list[756],sigma_out_list[757],sigma_out_list[758],sigma_out_list[759],sigma_out_list[760],sigma_out_list[761],sigma_out_list[762],sigma_out_list[763],sigma_out_list[764],sigma_out_list[765],sigma_out_list[766],sigma_out_list[767],sigma_out_list[768],sigma_out_list[769],sigma_out_list[770],sigma_out_list[771],sigma_out_list[772],sigma_out_list[773],sigma_out_list[774],sigma_out_list[775],sigma_out_list[776],sigma_out_list[777],sigma_out_list[778],sigma_out_list[779],sigma_out_list[780],sigma_out_list[781],sigma_out_list[782],sigma_out_list[783],sigma_out_list[784],sigma_out_list[785],sigma_out_list[786],sigma_out_list[787],sigma_out_list[788],sigma_out_list[789],sigma_out_list[790],sigma_out_list[791],sigma_out_list[792],sigma_out_list[793],sigma_out_list[794],sigma_out_list[795],sigma_out_list[796],sigma_out_list[797],sigma_out_list[798],sigma_out_list[799],sigma_out_list[800],sigma_out_list[801],sigma_out_list[802],sigma_out_list[803],sigma_out_list[804],sigma_out_list[805],sigma_out_list[806],sigma_out_list[807],sigma_out_list[808],sigma_out_list[809],sigma_out_list[810],sigma_out_list[811],sigma_out_list[812],sigma_out_list[813],sigma_out_list[814],sigma_out_list[815],sigma_out_list[816],sigma_out_list[817],sigma_out_list[818],sigma_out_list[819],sigma_out_list[820],sigma_out_list[821],sigma_out_list[822],sigma_out_list[823],sigma_out_list[824],sigma_out_list[825],sigma_out_list[826],sigma_out_list[827],sigma_out_list[828],sigma_out_list[829],sigma_out_list[830],sigma_out_list[831],sigma_out_list[832],sigma_out_list[833],sigma_out_list[834],sigma_out_list[835],sigma_out_list[836],sigma_out_list[837],sigma_out_list[838],sigma_out_list[839],sigma_out_list[840],sigma_out_list[841],sigma_out_list[842],sigma_out_list[843],sigma_out_list[844],sigma_out_list[845],sigma_out_list[846],sigma_out_list[847],sigma_out_list[848],sigma_out_list[849],sigma_out_list[850],sigma_out_list[851],sigma_out_list[852],sigma_out_list[853],sigma_out_list[854],sigma_out_list[855],sigma_out_list[856],sigma_out_list[857],sigma_out_list[858],sigma_out_list[859],sigma_out_list[860],sigma_out_list[861],sigma_out_list[862],sigma_out_list[863],sigma_out_list[864],sigma_out_list[865],sigma_out_list[866],sigma_out_list[867],sigma_out_list[868],sigma_out_list[869],sigma_out_list[870],sigma_out_list[871],sigma_out_list[872],sigma_out_list[873],sigma_out_list[874],sigma_out_list[875],sigma_out_list[876],sigma_out_list[877],sigma_out_list[878],sigma_out_list[879],sigma_out_list[880],sigma_out_list[881],sigma_out_list[882],sigma_out_list[883],sigma_out_list[884],sigma_out_list[885],sigma_out_list[886],sigma_out_list[887],sigma_out_list[888],sigma_out_list[889],sigma_out_list[890],sigma_out_list[891],sigma_out_list[892],sigma_out_list[893],sigma_out_list[894],sigma_out_list[895],sigma_out_list[896],sigma_out_list[897],sigma_out_list[898],sigma_out_list[899],sigma_out_list[900],sigma_out_list[901],sigma_out_list[902],sigma_out_list[903],sigma_out_list[904],sigma_out_list[905],sigma_out_list[906],sigma_out_list[907],sigma_out_list[908],sigma_out_list[909],sigma_out_list[910],sigma_out_list[911],sigma_out_list[912],sigma_out_list[913],sigma_out_list[914],sigma_out_list[915],sigma_out_list[916],sigma_out_list[917],sigma_out_list[918],sigma_out_list[919],sigma_out_list[920],sigma_out_list[921],sigma_out_list[922],sigma_out_list[923],sigma_out_list[924],sigma_out_list[925],sigma_out_list[926],sigma_out_list[927],sigma_out_list[928],sigma_out_list[929],sigma_out_list[930],sigma_out_list[931],sigma_out_list[932],sigma_out_list[933],sigma_out_list[934],sigma_out_list[935],sigma_out_list[936],sigma_out_list[937],sigma_out_list[938],sigma_out_list[939],sigma_out_list[940],sigma_out_list[941],sigma_out_list[942],sigma_out_list[943],sigma_out_list[944],sigma_out_list[945],sigma_out_list[946],sigma_out_list[947],sigma_out_list[948],sigma_out_list[949],sigma_out_list[950],sigma_out_list[951],sigma_out_list[952],sigma_out_list[953],sigma_out_list[954],sigma_out_list[955],sigma_out_list[956],sigma_out_list[957],sigma_out_list[958],sigma_out_list[959],sigma_out_list[960],sigma_out_list[961],sigma_out_list[962],sigma_out_list[963],sigma_out_list[964],sigma_out_list[965],sigma_out_list[966],sigma_out_list[967],sigma_out_list[968],sigma_out_list[969],sigma_out_list[970],sigma_out_list[971],sigma_out_list[972],sigma_out_list[973],sigma_out_list[974],sigma_out_list[975],sigma_out_list[976],sigma_out_list[977],sigma_out_list[978],sigma_out_list[979],sigma_out_list[980],sigma_out_list[981],sigma_out_list[982],sigma_out_list[983],sigma_out_list[984],sigma_out_list[985],sigma_out_list[986],sigma_out_list[987],sigma_out_list[988],sigma_out_list[989],sigma_out_list[990],sigma_out_list[991],sigma_out_list[992],sigma_out_list[993],sigma_out_list[994],sigma_out_list[995],sigma_out_list[996],sigma_out_list[997],sigma_out_list[998],sigma_out_list[999],sigma_out_list[1000],sigma_out_list[1001],sigma_out_list[1002],sigma_out_list[1003],sigma_out_list[1004],sigma_out_list[1005],sigma_out_list[1006],sigma_out_list[1007],sigma_out_list[1008],sigma_out_list[1009],sigma_out_list[1010],sigma_out_list[1011],sigma_out_list[1012],sigma_out_list[1013],sigma_out_list[1014],sigma_out_list[1015],sigma_out_list[1016],sigma_out_list[1017],sigma_out_list[1018],sigma_out_list[1019],sigma_out_list[1020],sigma_out_list[1021],sigma_out_list[1022],sigma_out_list[1023],sigma_out_list[1024],sigma_out_list[1025],sigma_out_list[1026],sigma_out_list[1027],sigma_out_list[1028],sigma_out_list[1029],sigma_out_list[1030],sigma_out_list[1031],sigma_out_list[1032],sigma_out_list[1033],sigma_out_list[1034],sigma_out_list[1035],sigma_out_list[1036],sigma_out_list[1037],sigma_out_list[1038],sigma_out_list[1039],sigma_out_list[1040],sigma_out_list[1041],sigma_out_list[1042],sigma_out_list[1043],sigma_out_list[1044],sigma_out_list[1045],sigma_out_list[1046],sigma_out_list[1047],sigma_out_list[1048],sigma_out_list[1049],sigma_out_list[1050],sigma_out_list[1051],sigma_out_list[1052],sigma_out_list[1053],sigma_out_list[1054],sigma_out_list[1055],sigma_out_list[1056],sigma_out_list[1057],sigma_out_list[1058],sigma_out_list[1059],sigma_out_list[1060],sigma_out_list[1061],sigma_out_list[1062],sigma_out_list[1063],sigma_out_list[1064],sigma_out_list[1065],sigma_out_list[1066],sigma_out_list[1067],sigma_out_list[1068],sigma_out_list[1069],sigma_out_list[1070],sigma_out_list[1071],sigma_out_list[1072],sigma_out_list[1073],sigma_out_list[1074],sigma_out_list[1075],sigma_out_list[1076],sigma_out_list[1077],sigma_out_list[1078],sigma_out_list[1079],sigma_out_list[1080],sigma_out_list[1081],sigma_out_list[1082],sigma_out_list[1083],sigma_out_list[1084],sigma_out_list[1085],sigma_out_list[1086],sigma_out_list[1087],sigma_out_list[1088],sigma_out_list[1089],sigma_out_list[1090],sigma_out_list[1091],sigma_out_list[1092],sigma_out_list[1093],sigma_out_list[1094],sigma_out_list[1095],sigma_out_list[1096],sigma_out_list[1097],sigma_out_list[1098],sigma_out_list[1099],sigma_out_list[1100],sigma_out_list[1101],sigma_out_list[1102],sigma_out_list[1103],sigma_out_list[1104],sigma_out_list[1105],sigma_out_list[1106],sigma_out_list[1107],sigma_out_list[1108],sigma_out_list[1109],sigma_out_list[1110],sigma_out_list[1111],sigma_out_list[1112],sigma_out_list[1113],sigma_out_list[1114],sigma_out_list[1115],sigma_out_list[1116],sigma_out_list[1117],sigma_out_list[1118],sigma_out_list[1119],sigma_out_list[1120],sigma_out_list[1121],sigma_out_list[1122],sigma_out_list[1123],sigma_out_list[1124],sigma_out_list[1125],sigma_out_list[1126],sigma_out_list[1127],sigma_out_list[1128],sigma_out_list[1129],sigma_out_list[1130],sigma_out_list[1131],sigma_out_list[1132],sigma_out_list[1133],sigma_out_list[1134],sigma_out_list[1135],sigma_out_list[1136],sigma_out_list[1137],sigma_out_list[1138],sigma_out_list[1139],sigma_out_list[1140],sigma_out_list[1141],sigma_out_list[1142],sigma_out_list[1143],sigma_out_list[1144],sigma_out_list[1145],sigma_out_list[1146],sigma_out_list[1147],sigma_out_list[1148],sigma_out_list[1149],sigma_out_list[1150],sigma_out_list[1151],sigma_out_list[1152],sigma_out_list[1153],sigma_out_list[1154],sigma_out_list[1155],sigma_out_list[1156],sigma_out_list[1157],sigma_out_list[1158],sigma_out_list[1159],sigma_out_list[1160],sigma_out_list[1161],sigma_out_list[1162],sigma_out_list[1163],sigma_out_list[1164],sigma_out_list[1165],sigma_out_list[1166],sigma_out_list[1167],sigma_out_list[1168],sigma_out_list[1169],sigma_out_list[1170],sigma_out_list[1171],sigma_out_list[1172],sigma_out_list[1173],sigma_out_list[1174],sigma_out_list[1175],sigma_out_list[1176],sigma_out_list[1177],sigma_out_list[1178],sigma_out_list[1179],sigma_out_list[1180],sigma_out_list[1181],sigma_out_list[1182],sigma_out_list[1183],sigma_out_list[1184],sigma_out_list[1185],sigma_out_list[1186],sigma_out_list[1187],sigma_out_list[1188],sigma_out_list[1189],sigma_out_list[1190],sigma_out_list[1191],sigma_out_list[1192],sigma_out_list[1193],sigma_out_list[1194],sigma_out_list[1195],sigma_out_list[1196],sigma_out_list[1197],sigma_out_list[1198],sigma_out_list[1199],sigma_out_list[1200],sigma_out_list[1201],sigma_out_list[1202],sigma_out_list[1203],sigma_out_list[1204],sigma_out_list[1205],sigma_out_list[1206],sigma_out_list[1207],sigma_out_list[1208],sigma_out_list[1209],sigma_out_list[1210],sigma_out_list[1211],sigma_out_list[1212],sigma_out_list[1213],sigma_out_list[1214],sigma_out_list[1215],sigma_out_list[1216],sigma_out_list[1217],sigma_out_list[1218],sigma_out_list[1219],sigma_out_list[1220],sigma_out_list[1221],sigma_out_list[1222],sigma_out_list[1223],sigma_out_list[1224],sigma_out_list[1225],sigma_out_list[1226],sigma_out_list[1227],sigma_out_list[1228],sigma_out_list[1229],sigma_out_list[1230],sigma_out_list[1231],sigma_out_list[1232],sigma_out_list[1233],sigma_out_list[1234],sigma_out_list[1235],sigma_out_list[1236],sigma_out_list[1237],sigma_out_list[1238],sigma_out_list[1239],sigma_out_list[1240],sigma_out_list[1241],sigma_out_list[1242],sigma_out_list[1243],sigma_out_list[1244],sigma_out_list[1245],sigma_out_list[1246],sigma_out_list[1247],sigma_out_list[1248],sigma_out_list[1249],sigma_out_list[1250],sigma_out_list[1251],sigma_out_list[1252],sigma_out_list[1253],sigma_out_list[1254],sigma_out_list[1255],sigma_out_list[1256],sigma_out_list[1257],sigma_out_list[1258],sigma_out_list[1259],sigma_out_list[1260],sigma_out_list[1261],sigma_out_list[1262],sigma_out_list[1263],sigma_out_list[1264],sigma_out_list[1265],sigma_out_list[1266],sigma_out_list[1267],sigma_out_list[1268],sigma_out_list[1269],sigma_out_list[1270],sigma_out_list[1271],sigma_out_list[1272],sigma_out_list[1273],sigma_out_list[1274],sigma_out_list[1275],sigma_out_list[1276],sigma_out_list[1277],sigma_out_list[1278],sigma_out_list[1279],sigma_out_list[1280],sigma_out_list[1281],sigma_out_list[1282],sigma_out_list[1283],sigma_out_list[1284],sigma_out_list[1285],sigma_out_list[1286],sigma_out_list[1287],sigma_out_list[1288],sigma_out_list[1289],sigma_out_list[1290],sigma_out_list[1291],sigma_out_list[1292],sigma_out_list[1293],sigma_out_list[1294],sigma_out_list[1295],sigma_out_list[1296],sigma_out_list[1297],sigma_out_list[1298],sigma_out_list[1299],sigma_out_list[1300],sigma_out_list[1301],sigma_out_list[1302],sigma_out_list[1303],sigma_out_list[1304],sigma_out_list[1305],sigma_out_list[1306],sigma_out_list[1307],sigma_out_list[1308],sigma_out_list[1309],sigma_out_list[1310],sigma_out_list[1311],sigma_out_list[1312],sigma_out_list[1313],sigma_out_list[1314],sigma_out_list[1315],sigma_out_list[1316],sigma_out_list[1317],sigma_out_list[1318],sigma_out_list[1319],sigma_out_list[1320],sigma_out_list[1321],sigma_out_list[1322],sigma_out_list[1323],sigma_out_list[1324],sigma_out_list[1325],sigma_out_list[1326],sigma_out_list[1327],sigma_out_list[1328],sigma_out_list[1329],sigma_out_list[1330],sigma_out_list[1331],sigma_out_list[1332],sigma_out_list[1333],sigma_out_list[1334],sigma_out_list[1335],sigma_out_list[1336],sigma_out_list[1337],sigma_out_list[1338],sigma_out_list[1339],sigma_out_list[1340],sigma_out_list[1341],sigma_out_list[1342],sigma_out_list[1343],sigma_out_list[1344],sigma_out_list[1345],sigma_out_list[1346],sigma_out_list[1347],sigma_out_list[1348],sigma_out_list[1349],sigma_out_list[1350],sigma_out_list[1351],sigma_out_list[1352],sigma_out_list[1353],sigma_out_list[1354],sigma_out_list[1355],sigma_out_list[1356],sigma_out_list[1357],sigma_out_list[1358],sigma_out_list[1359],sigma_out_list[1360],sigma_out_list[1361],sigma_out_list[1362],sigma_out_list[1363],sigma_out_list[1364],sigma_out_list[1365],sigma_out_list[1366],sigma_out_list[1367],sigma_out_list[1368],sigma_out_list[1369],sigma_out_list[1370],sigma_out_list[1371],sigma_out_list[1372],sigma_out_list[1373],sigma_out_list[1374],sigma_out_list[1375],sigma_out_list[1376],sigma_out_list[1377],sigma_out_list[1378],sigma_out_list[1379],sigma_out_list[1380],sigma_out_list[1381],sigma_out_list[1382],sigma_out_list[1383],sigma_out_list[1384],sigma_out_list[1385],sigma_out_list[1386],sigma_out_list[1387],sigma_out_list[1388],sigma_out_list[1389],sigma_out_list[1390],sigma_out_list[1391],sigma_out_list[1392],sigma_out_list[1393],sigma_out_list[1394],sigma_out_list[1395],sigma_out_list[1396],sigma_out_list[1397],sigma_out_list[1398],sigma_out_list[1399],sigma_out_list[1400],sigma_out_list[1401],sigma_out_list[1402],sigma_out_list[1403],sigma_out_list[1404],sigma_out_list[1405],sigma_out_list[1406],sigma_out_list[1407],sigma_out_list[1408],sigma_out_list[1409],sigma_out_list[1410],sigma_out_list[1411],sigma_out_list[1412],sigma_out_list[1413],sigma_out_list[1414],sigma_out_list[1415],sigma_out_list[1416],sigma_out_list[1417],sigma_out_list[1418],sigma_out_list[1419],sigma_out_list[1420],sigma_out_list[1421],sigma_out_list[1422],sigma_out_list[1423],sigma_out_list[1424],sigma_out_list[1425],sigma_out_list[1426],sigma_out_list[1427],sigma_out_list[1428],sigma_out_list[1429],sigma_out_list[1430],sigma_out_list[1431],sigma_out_list[1432],sigma_out_list[1433],sigma_out_list[1434],sigma_out_list[1435],sigma_out_list[1436],sigma_out_list[1437],sigma_out_list[1438],sigma_out_list[1439],sigma_out_list[1440],sigma_out_list[1441],sigma_out_list[1442],sigma_out_list[1443],sigma_out_list[1444],sigma_out_list[1445],sigma_out_list[1446],sigma_out_list[1447],sigma_out_list[1448],sigma_out_list[1449],sigma_out_list[1450],sigma_out_list[1451],sigma_out_list[1452],sigma_out_list[1453],sigma_out_list[1454],sigma_out_list[1455],sigma_out_list[1456],sigma_out_list[1457],sigma_out_list[1458],sigma_out_list[1459],sigma_out_list[1460],sigma_out_list[1461],sigma_out_list[1462],sigma_out_list[1463],sigma_out_list[1464],sigma_out_list[1465],sigma_out_list[1466],sigma_out_list[1467],sigma_out_list[1468],sigma_out_list[1469],sigma_out_list[1470],sigma_out_list[1471],sigma_out_list[1472],sigma_out_list[1473],sigma_out_list[1474],sigma_out_list[1475],sigma_out_list[1476],sigma_out_list[1477],sigma_out_list[1478],sigma_out_list[1479],sigma_out_list[1480],sigma_out_list[1481],sigma_out_list[1482],sigma_out_list[1483],sigma_out_list[1484],sigma_out_list[1485],sigma_out_list[1486],sigma_out_list[1487],sigma_out_list[1488],sigma_out_list[1489],sigma_out_list[1490],sigma_out_list[1491],sigma_out_list[1492],sigma_out_list[1493],sigma_out_list[1494],sigma_out_list[1495],sigma_out_list[1496],sigma_out_list[1497],sigma_out_list[1498],sigma_out_list[1499],sigma_out_list[1500],sigma_out_list[1501],sigma_out_list[1502],sigma_out_list[1503],sigma_out_list[1504],sigma_out_list[1505],sigma_out_list[1506],sigma_out_list[1507],sigma_out_list[1508],sigma_out_list[1509],sigma_out_list[1510],sigma_out_list[1511],sigma_out_list[1512],sigma_out_list[1513],sigma_out_list[1514],sigma_out_list[1515],sigma_out_list[1516],sigma_out_list[1517],sigma_out_list[1518],sigma_out_list[1519],sigma_out_list[1520],sigma_out_list[1521],sigma_out_list[1522],sigma_out_list[1523],sigma_out_list[1524],sigma_out_list[1525],sigma_out_list[1526],sigma_out_list[1527],sigma_out_list[1528],sigma_out_list[1529],sigma_out_list[1530],sigma_out_list[1531],sigma_out_list[1532],sigma_out_list[1533],sigma_out_list[1534],sigma_out_list[1535],sigma_out_list[1536],sigma_out_list[1537],sigma_out_list[1538],sigma_out_list[1539],sigma_out_list[1540],sigma_out_list[1541],sigma_out_list[1542],sigma_out_list[1543],sigma_out_list[1544],sigma_out_list[1545],sigma_out_list[1546],sigma_out_list[1547],sigma_out_list[1548],sigma_out_list[1549],sigma_out_list[1550],sigma_out_list[1551],sigma_out_list[1552],sigma_out_list[1553],sigma_out_list[1554],sigma_out_list[1555],sigma_out_list[1556],sigma_out_list[1557],sigma_out_list[1558],sigma_out_list[1559],sigma_out_list[1560],sigma_out_list[1561],sigma_out_list[1562],sigma_out_list[1563],sigma_out_list[1564],sigma_out_list[1565],sigma_out_list[1566],sigma_out_list[1567],sigma_out_list[1568],sigma_out_list[1569],sigma_out_list[1570],sigma_out_list[1571],sigma_out_list[1572],sigma_out_list[1573],sigma_out_list[1574],sigma_out_list[1575],sigma_out_list[1576],sigma_out_list[1577],sigma_out_list[1578],sigma_out_list[1579],sigma_out_list[1580],sigma_out_list[1581],sigma_out_list[1582],sigma_out_list[1583],sigma_out_list[1584],sigma_out_list[1585],sigma_out_list[1586],sigma_out_list[1587],sigma_out_list[1588],sigma_out_list[1589],sigma_out_list[1590],sigma_out_list[1591],sigma_out_list[1592],sigma_out_list[1593],sigma_out_list[1594],sigma_out_list[1595],sigma_out_list[1596],sigma_out_list[1597],sigma_out_list[1598],sigma_out_list[1599],sigma_out_list[1600],sigma_out_list[1601],sigma_out_list[1602],sigma_out_list[1603],sigma_out_list[1604],sigma_out_list[1605],sigma_out_list[1606],sigma_out_list[1607],sigma_out_list[1608],sigma_out_list[1609],sigma_out_list[1610],sigma_out_list[1611],sigma_out_list[1612],sigma_out_list[1613],sigma_out_list[1614],sigma_out_list[1615],sigma_out_list[1616],sigma_out_list[1617],sigma_out_list[1618],sigma_out_list[1619],sigma_out_list[1620],sigma_out_list[1621],sigma_out_list[1622],sigma_out_list[1623],sigma_out_list[1624],sigma_out_list[1625],sigma_out_list[1626],sigma_out_list[1627],sigma_out_list[1628],sigma_out_list[1629],sigma_out_list[1630],sigma_out_list[1631],sigma_out_list[1632],sigma_out_list[1633],sigma_out_list[1634],sigma_out_list[1635],sigma_out_list[1636],sigma_out_list[1637],sigma_out_list[1638],sigma_out_list[1639],sigma_out_list[1640],sigma_out_list[1641],sigma_out_list[1642],sigma_out_list[1643],sigma_out_list[1644],sigma_out_list[1645],sigma_out_list[1646],sigma_out_list[1647],sigma_out_list[1648],sigma_out_list[1649],sigma_out_list[1650],sigma_out_list[1651],sigma_out_list[1652],sigma_out_list[1653],sigma_out_list[1654],sigma_out_list[1655],sigma_out_list[1656],sigma_out_list[1657],sigma_out_list[1658],sigma_out_list[1659],sigma_out_list[1660],sigma_out_list[1661],sigma_out_list[1662],sigma_out_list[1663],sigma_out_list[1664],sigma_out_list[1665],sigma_out_list[1666],sigma_out_list[1667],sigma_out_list[1668],sigma_out_list[1669],sigma_out_list[1670],sigma_out_list[1671],sigma_out_list[1672],sigma_out_list[1673],sigma_out_list[1674],sigma_out_list[1675],sigma_out_list[1676],sigma_out_list[1677],sigma_out_list[1678],sigma_out_list[1679],sigma_out_list[1680],sigma_out_list[1681],sigma_out_list[1682],sigma_out_list[1683],sigma_out_list[1684],sigma_out_list[1685],sigma_out_list[1686],sigma_out_list[1687],sigma_out_list[1688],sigma_out_list[1689],sigma_out_list[1690],sigma_out_list[1691],sigma_out_list[1692],sigma_out_list[1693],sigma_out_list[1694],sigma_out_list[1695],sigma_out_list[1696],sigma_out_list[1697],sigma_out_list[1698],sigma_out_list[1699],sigma_out_list[1700],sigma_out_list[1701],sigma_out_list[1702],sigma_out_list[1703],sigma_out_list[1704],sigma_out_list[1705],sigma_out_list[1706],sigma_out_list[1707],sigma_out_list[1708],sigma_out_list[1709],sigma_out_list[1710],sigma_out_list[1711],sigma_out_list[1712],sigma_out_list[1713],sigma_out_list[1714],sigma_out_list[1715],sigma_out_list[1716],sigma_out_list[1717],sigma_out_list[1718],sigma_out_list[1719],sigma_out_list[1720],sigma_out_list[1721],sigma_out_list[1722],sigma_out_list[1723],sigma_out_list[1724],sigma_out_list[1725],sigma_out_list[1726],sigma_out_list[1727],sigma_out_list[1728],sigma_out_list[1729],sigma_out_list[1730],sigma_out_list[1731],sigma_out_list[1732],sigma_out_list[1733],sigma_out_list[1734],sigma_out_list[1735],sigma_out_list[1736],sigma_out_list[1737],sigma_out_list[1738],sigma_out_list[1739],sigma_out_list[1740],sigma_out_list[1741],sigma_out_list[1742],sigma_out_list[1743],sigma_out_list[1744],sigma_out_list[1745],sigma_out_list[1746],sigma_out_list[1747],sigma_out_list[1748],sigma_out_list[1749],sigma_out_list[1750],sigma_out_list[1751],sigma_out_list[1752],sigma_out_list[1753],sigma_out_list[1754],sigma_out_list[1755],sigma_out_list[1756],sigma_out_list[1757],sigma_out_list[1758],sigma_out_list[1759],sigma_out_list[1760],sigma_out_list[1761],sigma_out_list[1762],sigma_out_list[1763],sigma_out_list[1764],sigma_out_list[1765],sigma_out_list[1766],sigma_out_list[1767],sigma_out_list[1768],sigma_out_list[1769],sigma_out_list[1770],sigma_out_list[1771],sigma_out_list[1772],sigma_out_list[1773],sigma_out_list[1774],sigma_out_list[1775],sigma_out_list[1776],sigma_out_list[1777],sigma_out_list[1778],sigma_out_list[1779],sigma_out_list[1780],sigma_out_list[1781],sigma_out_list[1782],sigma_out_list[1783],sigma_out_list[1784],sigma_out_list[1785],sigma_out_list[1786],sigma_out_list[1787],sigma_out_list[1788],sigma_out_list[1789],sigma_out_list[1790],sigma_out_list[1791],sigma_out_list[1792],sigma_out_list[1793],sigma_out_list[1794],sigma_out_list[1795],sigma_out_list[1796],sigma_out_list[1797],sigma_out_list[1798],sigma_out_list[1799],sigma_out_list[1800],sigma_out_list[1801],sigma_out_list[1802],sigma_out_list[1803],sigma_out_list[1804],sigma_out_list[1805],sigma_out_list[1806],sigma_out_list[1807],sigma_out_list[1808],sigma_out_list[1809],sigma_out_list[1810],sigma_out_list[1811],sigma_out_list[1812],sigma_out_list[1813],sigma_out_list[1814],sigma_out_list[1815],sigma_out_list[1816],sigma_out_list[1817],sigma_out_list[1818],sigma_out_list[1819],sigma_out_list[1820],sigma_out_list[1821],sigma_out_list[1822],sigma_out_list[1823],sigma_out_list[1824],sigma_out_list[1825],sigma_out_list[1826],sigma_out_list[1827],sigma_out_list[1828],sigma_out_list[1829],sigma_out_list[1830],sigma_out_list[1831],sigma_out_list[1832],sigma_out_list[1833],sigma_out_list[1834],sigma_out_list[1835],sigma_out_list[1836],sigma_out_list[1837],sigma_out_list[1838],sigma_out_list[1839],sigma_out_list[1840],sigma_out_list[1841],sigma_out_list[1842],sigma_out_list[1843],sigma_out_list[1844],sigma_out_list[1845],sigma_out_list[1846],sigma_out_list[1847],sigma_out_list[1848],sigma_out_list[1849],sigma_out_list[1850],sigma_out_list[1851],sigma_out_list[1852],sigma_out_list[1853],sigma_out_list[1854],sigma_out_list[1855],sigma_out_list[1856],sigma_out_list[1857],sigma_out_list[1858],sigma_out_list[1859],sigma_out_list[1860],sigma_out_list[1861],sigma_out_list[1862],sigma_out_list[1863],sigma_out_list[1864],sigma_out_list[1865],sigma_out_list[1866],sigma_out_list[1867],sigma_out_list[1868],sigma_out_list[1869],sigma_out_list[1870],sigma_out_list[1871],sigma_out_list[1872],sigma_out_list[1873],sigma_out_list[1874],sigma_out_list[1875],sigma_out_list[1876],sigma_out_list[1877],sigma_out_list[1878],sigma_out_list[1879],sigma_out_list[1880],sigma_out_list[1881],sigma_out_list[1882],sigma_out_list[1883],sigma_out_list[1884],sigma_out_list[1885],sigma_out_list[1886],sigma_out_list[1887],sigma_out_list[1888],sigma_out_list[1889],sigma_out_list[1890],sigma_out_list[1891],sigma_out_list[1892],sigma_out_list[1893],sigma_out_list[1894],sigma_out_list[1895],sigma_out_list[1896],sigma_out_list[1897],sigma_out_list[1898],sigma_out_list[1899],sigma_out_list[1900],sigma_out_list[1901],sigma_out_list[1902],sigma_out_list[1903],sigma_out_list[1904],sigma_out_list[1905],sigma_out_list[1906],sigma_out_list[1907],sigma_out_list[1908],sigma_out_list[1909],sigma_out_list[1910],sigma_out_list[1911],sigma_out_list[1912],sigma_out_list[1913],sigma_out_list[1914],sigma_out_list[1915],sigma_out_list[1916],sigma_out_list[1917],sigma_out_list[1918],sigma_out_list[1919],sigma_out_list[1920],sigma_out_list[1921],sigma_out_list[1922],sigma_out_list[1923],sigma_out_list[1924],sigma_out_list[1925],sigma_out_list[1926],sigma_out_list[1927],sigma_out_list[1928],sigma_out_list[1929],sigma_out_list[1930],sigma_out_list[1931],sigma_out_list[1932],sigma_out_list[1933],sigma_out_list[1934],sigma_out_list[1935],sigma_out_list[1936],sigma_out_list[1937],sigma_out_list[1938],sigma_out_list[1939],sigma_out_list[1940],sigma_out_list[1941],sigma_out_list[1942],sigma_out_list[1943],sigma_out_list[1944],sigma_out_list[1945],sigma_out_list[1946],sigma_out_list[1947],sigma_out_list[1948],sigma_out_list[1949],sigma_out_list[1950],sigma_out_list[1951],sigma_out_list[1952],sigma_out_list[1953],sigma_out_list[1954],sigma_out_list[1955],sigma_out_list[1956],sigma_out_list[1957],sigma_out_list[1958],sigma_out_list[1959],sigma_out_list[1960],sigma_out_list[1961],sigma_out_list[1962],sigma_out_list[1963],sigma_out_list[1964],sigma_out_list[1965],sigma_out_list[1966],sigma_out_list[1967],sigma_out_list[1968],sigma_out_list[1969],sigma_out_list[1970],sigma_out_list[1971],sigma_out_list[1972],sigma_out_list[1973],sigma_out_list[1974],sigma_out_list[1975],sigma_out_list[1976],sigma_out_list[1977],sigma_out_list[1978],sigma_out_list[1979],sigma_out_list[1980],sigma_out_list[1981],sigma_out_list[1982],sigma_out_list[1983],sigma_out_list[1984],sigma_out_list[1985],sigma_out_list[1986],sigma_out_list[1987],sigma_out_list[1988],sigma_out_list[1989],sigma_out_list[1990],sigma_out_list[1991],sigma_out_list[1992],sigma_out_list[1993],sigma_out_list[1994],sigma_out_list[1995],sigma_out_list[1996],sigma_out_list[1997],sigma_out_list[1998],sigma_out_list[1999],sigma_out_list[2000],sigma_out_list[2001],sigma_out_list[2002],sigma_out_list[2003],sigma_out_list[2004],sigma_out_list[2005],sigma_out_list[2006],sigma_out_list[2007],sigma_out_list[2008],sigma_out_list[2009],sigma_out_list[2010],sigma_out_list[2011],sigma_out_list[2012],sigma_out_list[2013],sigma_out_list[2014],sigma_out_list[2015],sigma_out_list[2016],sigma_out_list[2017],sigma_out_list[2018],sigma_out_list[2019],sigma_out_list[2020],sigma_out_list[2021],sigma_out_list[2022],sigma_out_list[2023],sigma_out_list[2024],sigma_out_list[2025],sigma_out_list[2026],sigma_out_list[2027],sigma_out_list[2028],sigma_out_list[2029],sigma_out_list[2030],sigma_out_list[2031],sigma_out_list[2032],sigma_out_list[2033],sigma_out_list[2034],sigma_out_list[2035],sigma_out_list[2036],sigma_out_list[2037],sigma_out_list[2038],sigma_out_list[2039],sigma_out_list[2040],sigma_out_list[2041],sigma_out_list[2042],sigma_out_list[2043],sigma_out_list[2044],sigma_out_list[2045],sigma_out_list[2046],sigma_out_list[2047],sigma_out_list[2048],sigma_out_list[2049],sigma_out_list[2050],sigma_out_list[2051],sigma_out_list[2052],sigma_out_list[2053],sigma_out_list[2054],sigma_out_list[2055],sigma_out_list[2056],sigma_out_list[2057],sigma_out_list[2058],sigma_out_list[2059],sigma_out_list[2060],sigma_out_list[2061],sigma_out_list[2062],sigma_out_list[2063],sigma_out_list[2064],sigma_out_list[2065],sigma_out_list[2066],sigma_out_list[2067],sigma_out_list[2068],sigma_out_list[2069],sigma_out_list[2070],sigma_out_list[2071],sigma_out_list[2072],sigma_out_list[2073],sigma_out_list[2074],sigma_out_list[2075],sigma_out_list[2076],sigma_out_list[2077],sigma_out_list[2078],sigma_out_list[2079],sigma_out_list[2080],sigma_out_list[2081],sigma_out_list[2082],sigma_out_list[2083],sigma_out_list[2084],sigma_out_list[2085],sigma_out_list[2086],sigma_out_list[2087],sigma_out_list[2088],sigma_out_list[2089],sigma_out_list[2090],sigma_out_list[2091],sigma_out_list[2092],sigma_out_list[2093],sigma_out_list[2094],sigma_out_list[2095],sigma_out_list[2096],sigma_out_list[2097],sigma_out_list[2098],sigma_out_list[2099],sigma_out_list[2100],sigma_out_list[2101],sigma_out_list[2102],sigma_out_list[2103],sigma_out_list[2104],sigma_out_list[2105],sigma_out_list[2106],sigma_out_list[2107],sigma_out_list[2108],sigma_out_list[2109],sigma_out_list[2110],sigma_out_list[2111],sigma_out_list[2112],sigma_out_list[2113],sigma_out_list[2114],sigma_out_list[2115],sigma_out_list[2116],sigma_out_list[2117],sigma_out_list[2118],sigma_out_list[2119],sigma_out_list[2120],sigma_out_list[2121],sigma_out_list[2122],sigma_out_list[2123],sigma_out_list[2124],sigma_out_list[2125],sigma_out_list[2126],sigma_out_list[2127],sigma_out_list[2128],sigma_out_list[2129],sigma_out_list[2130],sigma_out_list[2131],sigma_out_list[2132],sigma_out_list[2133],sigma_out_list[2134],sigma_out_list[2135],sigma_out_list[2136],sigma_out_list[2137],sigma_out_list[2138],sigma_out_list[2139],sigma_out_list[2140],sigma_out_list[2141],sigma_out_list[2142],sigma_out_list[2143],sigma_out_list[2144],sigma_out_list[2145],sigma_out_list[2146],sigma_out_list[2147],sigma_out_list[2148],sigma_out_list[2149],sigma_out_list[2150],sigma_out_list[2151],sigma_out_list[2152],sigma_out_list[2153],sigma_out_list[2154],sigma_out_list[2155],sigma_out_list[2156],sigma_out_list[2157],sigma_out_list[2158],sigma_out_list[2159],sigma_out_list[2160],sigma_out_list[2161],sigma_out_list[2162],sigma_out_list[2163],sigma_out_list[2164],sigma_out_list[2165],sigma_out_list[2166],sigma_out_list[2167],sigma_out_list[2168],sigma_out_list[2169],sigma_out_list[2170],sigma_out_list[2171],sigma_out_list[2172],sigma_out_list[2173],sigma_out_list[2174],sigma_out_list[2175],sigma_out_list[2176],sigma_out_list[2177],sigma_out_list[2178],sigma_out_list[2179],sigma_out_list[2180],sigma_out_list[2181],sigma_out_list[2182],sigma_out_list[2183],sigma_out_list[2184],sigma_out_list[2185],sigma_out_list[2186],sigma_out_list[2187],sigma_out_list[2188],sigma_out_list[2189],sigma_out_list[2190],sigma_out_list[2191],sigma_out_list[2192],sigma_out_list[2193],sigma_out_list[2194],sigma_out_list[2195],sigma_out_list[2196],sigma_out_list[2197],sigma_out_list[2198],sigma_out_list[2199],sigma_out_list[2200],sigma_out_list[2201],sigma_out_list[2202],sigma_out_list[2203],sigma_out_list[2204],sigma_out_list[2205],sigma_out_list[2206],sigma_out_list[2207],sigma_out_list[2208],sigma_out_list[2209],sigma_out_list[2210],sigma_out_list[2211],sigma_out_list[2212],sigma_out_list[2213],sigma_out_list[2214],sigma_out_list[2215],sigma_out_list[2216],sigma_out_list[2217],sigma_out_list[2218],sigma_out_list[2219],sigma_out_list[2220],sigma_out_list[2221],sigma_out_list[2222],sigma_out_list[2223],sigma_out_list[2224],sigma_out_list[2225],sigma_out_list[2226],sigma_out_list[2227],sigma_out_list[2228],sigma_out_list[2229],sigma_out_list[2230],sigma_out_list[2231],sigma_out_list[2232],sigma_out_list[2233],sigma_out_list[2234],sigma_out_list[2235],sigma_out_list[2236],sigma_out_list[2237],sigma_out_list[2238],sigma_out_list[2239],sigma_out_list[2240],sigma_out_list[2241],sigma_out_list[2242],sigma_out_list[2243],sigma_out_list[2244],sigma_out_list[2245],sigma_out_list[2246],sigma_out_list[2247],sigma_out_list[2248],sigma_out_list[2249],sigma_out_list[2250],sigma_out_list[2251],sigma_out_list[2252],sigma_out_list[2253],sigma_out_list[2254],sigma_out_list[2255],sigma_out_list[2256],sigma_out_list[2257],sigma_out_list[2258],sigma_out_list[2259],sigma_out_list[2260],sigma_out_list[2261],sigma_out_list[2262],sigma_out_list[2263],sigma_out_list[2264],sigma_out_list[2265],sigma_out_list[2266],sigma_out_list[2267],sigma_out_list[2268],sigma_out_list[2269],sigma_out_list[2270],sigma_out_list[2271],sigma_out_list[2272],sigma_out_list[2273],sigma_out_list[2274],sigma_out_list[2275],sigma_out_list[2276],sigma_out_list[2277],sigma_out_list[2278],sigma_out_list[2279],sigma_out_list[2280],sigma_out_list[2281],sigma_out_list[2282],sigma_out_list[2283],sigma_out_list[2284],sigma_out_list[2285],sigma_out_list[2286],sigma_out_list[2287],sigma_out_list[2288],sigma_out_list[2289],sigma_out_list[2290],sigma_out_list[2291],sigma_out_list[2292],sigma_out_list[2293],sigma_out_list[2294],sigma_out_list[2295],sigma_out_list[2296],sigma_out_list[2297],sigma_out_list[2298],sigma_out_list[2299],sigma_out_list[2300],sigma_out_list[2301],sigma_out_list[2302],sigma_out_list[2303],sigma_out_list[2304],sigma_out_list[2305],sigma_out_list[2306],sigma_out_list[2307],sigma_out_list[2308],sigma_out_list[2309],sigma_out_list[2310],sigma_out_list[2311],sigma_out_list[2312],sigma_out_list[2313],sigma_out_list[2314],sigma_out_list[2315],sigma_out_list[2316],sigma_out_list[2317],sigma_out_list[2318],sigma_out_list[2319],sigma_out_list[2320],sigma_out_list[2321],sigma_out_list[2322],sigma_out_list[2323],sigma_out_list[2324],sigma_out_list[2325],sigma_out_list[2326],sigma_out_list[2327],sigma_out_list[2328],sigma_out_list[2329],sigma_out_list[2330],sigma_out_list[2331],sigma_out_list[2332],sigma_out_list[2333],sigma_out_list[2334],sigma_out_list[2335],sigma_out_list[2336],sigma_out_list[2337],sigma_out_list[2338],sigma_out_list[2339],sigma_out_list[2340],sigma_out_list[2341],sigma_out_list[2342],sigma_out_list[2343],sigma_out_list[2344],sigma_out_list[2345],sigma_out_list[2346],sigma_out_list[2347],sigma_out_list[2348],sigma_out_list[2349],sigma_out_list[2350],sigma_out_list[2351],sigma_out_list[2352],sigma_out_list[2353],sigma_out_list[2354],sigma_out_list[2355],sigma_out_list[2356],sigma_out_list[2357],sigma_out_list[2358],sigma_out_list[2359],sigma_out_list[2360],sigma_out_list[2361],sigma_out_list[2362],sigma_out_list[2363],sigma_out_list[2364],sigma_out_list[2365],sigma_out_list[2366],sigma_out_list[2367],sigma_out_list[2368],sigma_out_list[2369],sigma_out_list[2370],sigma_out_list[2371],sigma_out_list[2372],sigma_out_list[2373],sigma_out_list[2374],sigma_out_list[2375],sigma_out_list[2376],sigma_out_list[2377],sigma_out_list[2378],sigma_out_list[2379],sigma_out_list[2380],sigma_out_list[2381],sigma_out_list[2382],sigma_out_list[2383],sigma_out_list[2384],sigma_out_list[2385],sigma_out_list[2386],sigma_out_list[2387],sigma_out_list[2388],sigma_out_list[2389],sigma_out_list[2390],sigma_out_list[2391],sigma_out_list[2392],sigma_out_list[2393],sigma_out_list[2394],sigma_out_list[2395],sigma_out_list[2396],sigma_out_list[2397],sigma_out_list[2398],sigma_out_list[2399],sigma_out_list[2400],sigma_out_list[2401],sigma_out_list[2402],sigma_out_list[2403],sigma_out_list[2404],sigma_out_list[2405],sigma_out_list[2406],sigma_out_list[2407],sigma_out_list[2408],sigma_out_list[2409],sigma_out_list[2410],sigma_out_list[2411],sigma_out_list[2412],sigma_out_list[2413],sigma_out_list[2414],sigma_out_list[2415],sigma_out_list[2416],sigma_out_list[2417],sigma_out_list[2418],sigma_out_list[2419],sigma_out_list[2420],sigma_out_list[2421],sigma_out_list[2422],sigma_out_list[2423],sigma_out_list[2424],sigma_out_list[2425],sigma_out_list[2426],sigma_out_list[2427],sigma_out_list[2428],sigma_out_list[2429],sigma_out_list[2430],sigma_out_list[2431],sigma_out_list[2432],sigma_out_list[2433],sigma_out_list[2434],sigma_out_list[2435],sigma_out_list[2436],sigma_out_list[2437],sigma_out_list[2438],sigma_out_list[2439],sigma_out_list[2440],sigma_out_list[2441],sigma_out_list[2442],sigma_out_list[2443],sigma_out_list[2444],sigma_out_list[2445],sigma_out_list[2446],sigma_out_list[2447]}=sigma_out;



always @(posedge sys_clk or negedge sys_rst_n)begin
	if(!sys_rst_n)begin
		counter<=0;
		wea<=0;
		w_ram_from_sign_end<=0;
		state<=0;
	end
	else begin
	    if(~w_ram_from_sign_start) begin
	       w_ram_from_sign_end<=0;
	    end
	    if(w_ram_from_sign_start==1&&state==0&&w_ram_from_sign_end==0)begin
			data<=sigma_out_list[counter];
			wea<=1;
			state<=1;
		end
		else if(state==1) begin
			state<=2;
		end
		else if(state==2) begin
			counter<=counter+1;
			wea<=0;
			if(counter==full_number-1) begin
				state<=3;
			end
			else begin
				state<=0;
			end
		end
		else if(state==3) begin
		    wea<=0;
			counter<=0;
			w_ram_from_sign_end<=1;
			state<=0;
		end
	end
end

endmodule

