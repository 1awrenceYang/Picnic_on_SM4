/*
    input clk,
    input reset,
    input[0:3] mode,
    input[0:2*1088-1] h1InSeedSet,
    input Hstart,
    input[0:9] groupNum,
    output [0:511] hashValue,
    output reg en_end
*/

module seed_tree(
    input clk,
    input reset,
    //input root_seed,
    //input salt
    input tree_start,
    output reg [256*602-1:0] iseed,
    output reg tree_set_end
    );
    wire [0:255] salt=0;
    reg [2*1088-1:0] h1InSeedSet [300:0];
    wire t=1;
    wire j=1;
    wire [573+1088:0]padding=0;
    reg [300:0] Hstart;
    reg [300:0] restart;
    wire [511:0] hashValue[300:0];
    wire [300:0] en_end;
    wire [9:0] groupNum=2;
    reg[4:0] state; 
    reg[9:0] counter;
    wire [0:300] start_marsk[0:9];
    assign start_marsk[0] = 1;
    assign start_marsk[1] = 301'h3;
    assign start_marsk[2] = 301'hf;
    assign start_marsk[3] = 301'hff;
    assign start_marsk[4] = 301'hffff;
    assign start_marsk[5] = 301'hffffffff;
    assign start_marsk[6] = 301'hffffffffffffffff;
    assign start_marsk[7] = 301'hffffffffffffffffffffffffffffffff;
    assign start_marsk[8] = 301'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
    assign start_marsk[9] = 301'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;

    always @(posedge clk or negedge reset) begin
        if(~reset) begin
            counter <= 0;
            state<=0;
            tree_set_end<=0;
        end
        else begin
            if(state==0) begin
                if(tree_start) begin
                    tree_set_end<=0;
                    Hstart<=start_marsk[counter];
                    restart<=0;
                    state<=1;
                    if(counter==0)begin
                        //h1InSeedSet[0]={root_seed,salt,t,j,padding};
                        h1InSeedSet[0]<=0;
                    end
                end
                
            end
            if(state==1) begin
                if(en_end==start_marsk[counter]) begin
                        counter<=counter+1;
                        restart<=Hstart;
                        if(en_end == start_marsk[9]) begin
                            state<=2;
                        end
                        else begin
                            state<=0;
                        end
                        h1InSeedSet[0]<={hashValue[0][511:256],salt,t,j,padding};
                        h1InSeedSet[1]<={hashValue[0][255:0],salt,t,j,padding};
                        h1InSeedSet[2]<={hashValue[1][511:256],salt,t,j,padding};
                        h1InSeedSet[3]<={hashValue[1][255:0],salt,t,j,padding};
                        h1InSeedSet[4]<={hashValue[2][511:256],salt,t,j,padding};
                        h1InSeedSet[5]<={hashValue[2][255:0],salt,t,j,padding};
                        h1InSeedSet[6]<={hashValue[3][511:256],salt,t,j,padding};
                        h1InSeedSet[7]<={hashValue[3][255:0],salt,t,j,padding};
                        h1InSeedSet[8]<={hashValue[4][511:256],salt,t,j,padding};
                        h1InSeedSet[9]<={hashValue[4][255:0],salt,t,j,padding};
                        h1InSeedSet[10]<={hashValue[5][511:256],salt,t,j,padding};
                        h1InSeedSet[11]<={hashValue[5][255:0],salt,t,j,padding};
                        h1InSeedSet[12]<={hashValue[6][511:256],salt,t,j,padding};
                        h1InSeedSet[13]<={hashValue[6][255:0],salt,t,j,padding};
                        h1InSeedSet[14]<={hashValue[7][511:256],salt,t,j,padding};
                        h1InSeedSet[15]<={hashValue[7][255:0],salt,t,j,padding};
                        h1InSeedSet[16]<={hashValue[8][511:256],salt,t,j,padding};
                        h1InSeedSet[17]<={hashValue[8][255:0],salt,t,j,padding};
                        h1InSeedSet[18]<={hashValue[9][511:256],salt,t,j,padding};
                        h1InSeedSet[19]<={hashValue[9][255:0],salt,t,j,padding};
                        h1InSeedSet[20]<={hashValue[10][511:256],salt,t,j,padding};
                        h1InSeedSet[21]<={hashValue[10][255:0],salt,t,j,padding};
                        h1InSeedSet[22]<={hashValue[11][511:256],salt,t,j,padding};
                        h1InSeedSet[23]<={hashValue[11][255:0],salt,t,j,padding};
                        h1InSeedSet[24]<={hashValue[12][511:256],salt,t,j,padding};
                        h1InSeedSet[25]<={hashValue[12][255:0],salt,t,j,padding};
                        h1InSeedSet[26]<={hashValue[13][511:256],salt,t,j,padding};
                        h1InSeedSet[27]<={hashValue[13][255:0],salt,t,j,padding};
                        h1InSeedSet[28]<={hashValue[14][511:256],salt,t,j,padding};
                        h1InSeedSet[29]<={hashValue[14][255:0],salt,t,j,padding};
                        h1InSeedSet[30]<={hashValue[15][511:256],salt,t,j,padding};
                        h1InSeedSet[31]<={hashValue[15][255:0],salt,t,j,padding};
                        h1InSeedSet[32]<={hashValue[16][511:256],salt,t,j,padding};
                        h1InSeedSet[33]<={hashValue[16][255:0],salt,t,j,padding};
                        h1InSeedSet[34]<={hashValue[17][511:256],salt,t,j,padding};
                        h1InSeedSet[35]<={hashValue[17][255:0],salt,t,j,padding};
                        h1InSeedSet[36]<={hashValue[18][511:256],salt,t,j,padding};
                        h1InSeedSet[37]<={hashValue[18][255:0],salt,t,j,padding};
                        h1InSeedSet[38]<={hashValue[19][511:256],salt,t,j,padding};
                        h1InSeedSet[39]<={hashValue[19][255:0],salt,t,j,padding};
                        h1InSeedSet[40]<={hashValue[20][511:256],salt,t,j,padding};
                        h1InSeedSet[41]<={hashValue[20][255:0],salt,t,j,padding};
                        h1InSeedSet[42]<={hashValue[21][511:256],salt,t,j,padding};
                        h1InSeedSet[43]<={hashValue[21][255:0],salt,t,j,padding};
                        h1InSeedSet[44]<={hashValue[22][511:256],salt,t,j,padding};
                        h1InSeedSet[45]<={hashValue[22][255:0],salt,t,j,padding};
                        h1InSeedSet[46]<={hashValue[23][511:256],salt,t,j,padding};
                        h1InSeedSet[47]<={hashValue[23][255:0],salt,t,j,padding};
                        h1InSeedSet[48]<={hashValue[24][511:256],salt,t,j,padding};
                        h1InSeedSet[49]<={hashValue[24][255:0],salt,t,j,padding};
                        h1InSeedSet[50]<={hashValue[25][511:256],salt,t,j,padding};
                        h1InSeedSet[51]<={hashValue[25][255:0],salt,t,j,padding};
                        h1InSeedSet[52]<={hashValue[26][511:256],salt,t,j,padding};
                        h1InSeedSet[53]<={hashValue[26][255:0],salt,t,j,padding};
                        h1InSeedSet[54]<={hashValue[27][511:256],salt,t,j,padding};
                        h1InSeedSet[55]<={hashValue[27][255:0],salt,t,j,padding};
                        h1InSeedSet[56]<={hashValue[28][511:256],salt,t,j,padding};
                        h1InSeedSet[57]<={hashValue[28][255:0],salt,t,j,padding};
                        h1InSeedSet[58]<={hashValue[29][511:256],salt,t,j,padding};
                        h1InSeedSet[59]<={hashValue[29][255:0],salt,t,j,padding};
                        h1InSeedSet[60]<={hashValue[30][511:256],salt,t,j,padding};
                        h1InSeedSet[61]<={hashValue[30][255:0],salt,t,j,padding};
                        h1InSeedSet[62]<={hashValue[31][511:256],salt,t,j,padding};
                        h1InSeedSet[63]<={hashValue[31][255:0],salt,t,j,padding};
                        h1InSeedSet[64]<={hashValue[32][511:256],salt,t,j,padding};
                        h1InSeedSet[65]<={hashValue[32][255:0],salt,t,j,padding};
                        h1InSeedSet[66]<={hashValue[33][511:256],salt,t,j,padding};
                        h1InSeedSet[67]<={hashValue[33][255:0],salt,t,j,padding};
                        h1InSeedSet[68]<={hashValue[34][511:256],salt,t,j,padding};
                        h1InSeedSet[69]<={hashValue[34][255:0],salt,t,j,padding};
                        h1InSeedSet[70]<={hashValue[35][511:256],salt,t,j,padding};
                        h1InSeedSet[71]<={hashValue[35][255:0],salt,t,j,padding};
                        h1InSeedSet[72]<={hashValue[36][511:256],salt,t,j,padding};
                        h1InSeedSet[73]<={hashValue[36][255:0],salt,t,j,padding};
                        h1InSeedSet[74]<={hashValue[37][511:256],salt,t,j,padding};
                        h1InSeedSet[75]<={hashValue[37][255:0],salt,t,j,padding};
                        h1InSeedSet[76]<={hashValue[38][511:256],salt,t,j,padding};
                        h1InSeedSet[77]<={hashValue[38][255:0],salt,t,j,padding};
                        h1InSeedSet[78]<={hashValue[39][511:256],salt,t,j,padding};
                        h1InSeedSet[79]<={hashValue[39][255:0],salt,t,j,padding};
                        h1InSeedSet[80]<={hashValue[40][511:256],salt,t,j,padding};
                        h1InSeedSet[81]<={hashValue[40][255:0],salt,t,j,padding};
                        h1InSeedSet[82]<={hashValue[41][511:256],salt,t,j,padding};
                        h1InSeedSet[83]<={hashValue[41][255:0],salt,t,j,padding};
                        h1InSeedSet[84]<={hashValue[42][511:256],salt,t,j,padding};
                        h1InSeedSet[85]<={hashValue[42][255:0],salt,t,j,padding};
                        h1InSeedSet[86]<={hashValue[43][511:256],salt,t,j,padding};
                        h1InSeedSet[87]<={hashValue[43][255:0],salt,t,j,padding};
                        h1InSeedSet[88]<={hashValue[44][511:256],salt,t,j,padding};
                        h1InSeedSet[89]<={hashValue[44][255:0],salt,t,j,padding};
                        h1InSeedSet[90]<={hashValue[45][511:256],salt,t,j,padding};
                        h1InSeedSet[91]<={hashValue[45][255:0],salt,t,j,padding};
                        h1InSeedSet[92]<={hashValue[46][511:256],salt,t,j,padding};
                        h1InSeedSet[93]<={hashValue[46][255:0],salt,t,j,padding};
                        h1InSeedSet[94]<={hashValue[47][511:256],salt,t,j,padding};
                        h1InSeedSet[95]<={hashValue[47][255:0],salt,t,j,padding};
                        h1InSeedSet[96]<={hashValue[48][511:256],salt,t,j,padding};
                        h1InSeedSet[97]<={hashValue[48][255:0],salt,t,j,padding};
                        h1InSeedSet[98]<={hashValue[49][511:256],salt,t,j,padding};
                        h1InSeedSet[99]<={hashValue[49][255:0],salt,t,j,padding};
                        h1InSeedSet[100]<={hashValue[50][511:256],salt,t,j,padding};
                        h1InSeedSet[101]<={hashValue[50][255:0],salt,t,j,padding};
                        h1InSeedSet[102]<={hashValue[51][511:256],salt,t,j,padding};
                        h1InSeedSet[103]<={hashValue[51][255:0],salt,t,j,padding};
                        h1InSeedSet[104]<={hashValue[52][511:256],salt,t,j,padding};
                        h1InSeedSet[105]<={hashValue[52][255:0],salt,t,j,padding};
                        h1InSeedSet[106]<={hashValue[53][511:256],salt,t,j,padding};
                        h1InSeedSet[107]<={hashValue[53][255:0],salt,t,j,padding};
                        h1InSeedSet[108]<={hashValue[54][511:256],salt,t,j,padding};
                        h1InSeedSet[109]<={hashValue[54][255:0],salt,t,j,padding};
                        h1InSeedSet[110]<={hashValue[55][511:256],salt,t,j,padding};
                        h1InSeedSet[111]<={hashValue[55][255:0],salt,t,j,padding};
                        h1InSeedSet[112]<={hashValue[56][511:256],salt,t,j,padding};
                        h1InSeedSet[113]<={hashValue[56][255:0],salt,t,j,padding};
                        h1InSeedSet[114]<={hashValue[57][511:256],salt,t,j,padding};
                        h1InSeedSet[115]<={hashValue[57][255:0],salt,t,j,padding};
                        h1InSeedSet[116]<={hashValue[58][511:256],salt,t,j,padding};
                        h1InSeedSet[117]<={hashValue[58][255:0],salt,t,j,padding};
                        h1InSeedSet[118]<={hashValue[59][511:256],salt,t,j,padding};
                        h1InSeedSet[119]<={hashValue[59][255:0],salt,t,j,padding};
                        h1InSeedSet[120]<={hashValue[60][511:256],salt,t,j,padding};
                        h1InSeedSet[121]<={hashValue[60][255:0],salt,t,j,padding};
                        h1InSeedSet[122]<={hashValue[61][511:256],salt,t,j,padding};
                        h1InSeedSet[123]<={hashValue[61][255:0],salt,t,j,padding};
                        h1InSeedSet[124]<={hashValue[62][511:256],salt,t,j,padding};
                        h1InSeedSet[125]<={hashValue[62][255:0],salt,t,j,padding};
                        h1InSeedSet[126]<={hashValue[63][511:256],salt,t,j,padding};
                        h1InSeedSet[127]<={hashValue[63][255:0],salt,t,j,padding};
                        h1InSeedSet[128]<={hashValue[64][511:256],salt,t,j,padding};
                        h1InSeedSet[129]<={hashValue[64][255:0],salt,t,j,padding};
                        h1InSeedSet[130]<={hashValue[65][511:256],salt,t,j,padding};
                        h1InSeedSet[131]<={hashValue[65][255:0],salt,t,j,padding};
                        h1InSeedSet[132]<={hashValue[66][511:256],salt,t,j,padding};
                        h1InSeedSet[133]<={hashValue[66][255:0],salt,t,j,padding};
                        h1InSeedSet[134]<={hashValue[67][511:256],salt,t,j,padding};
                        h1InSeedSet[135]<={hashValue[67][255:0],salt,t,j,padding};
                        h1InSeedSet[136]<={hashValue[68][511:256],salt,t,j,padding};
                        h1InSeedSet[137]<={hashValue[68][255:0],salt,t,j,padding};
                        h1InSeedSet[138]<={hashValue[69][511:256],salt,t,j,padding};
                        h1InSeedSet[139]<={hashValue[69][255:0],salt,t,j,padding};
                        h1InSeedSet[140]<={hashValue[70][511:256],salt,t,j,padding};
                        h1InSeedSet[141]<={hashValue[70][255:0],salt,t,j,padding};
                        h1InSeedSet[142]<={hashValue[71][511:256],salt,t,j,padding};
                        h1InSeedSet[143]<={hashValue[71][255:0],salt,t,j,padding};
                        h1InSeedSet[144]<={hashValue[72][511:256],salt,t,j,padding};
                        h1InSeedSet[145]<={hashValue[72][255:0],salt,t,j,padding};
                        h1InSeedSet[146]<={hashValue[73][511:256],salt,t,j,padding};
                        h1InSeedSet[147]<={hashValue[73][255:0],salt,t,j,padding};
                        h1InSeedSet[148]<={hashValue[74][511:256],salt,t,j,padding};
                        h1InSeedSet[149]<={hashValue[74][255:0],salt,t,j,padding};
                        h1InSeedSet[150]<={hashValue[75][511:256],salt,t,j,padding};
                        h1InSeedSet[151]<={hashValue[75][255:0],salt,t,j,padding};
                        h1InSeedSet[152]<={hashValue[76][511:256],salt,t,j,padding};
                        h1InSeedSet[153]<={hashValue[76][255:0],salt,t,j,padding};
                        h1InSeedSet[154]<={hashValue[77][511:256],salt,t,j,padding};
                        h1InSeedSet[155]<={hashValue[77][255:0],salt,t,j,padding};
                        h1InSeedSet[156]<={hashValue[78][511:256],salt,t,j,padding};
                        h1InSeedSet[157]<={hashValue[78][255:0],salt,t,j,padding};
                        h1InSeedSet[158]<={hashValue[79][511:256],salt,t,j,padding};
                        h1InSeedSet[159]<={hashValue[79][255:0],salt,t,j,padding};
                        h1InSeedSet[160]<={hashValue[80][511:256],salt,t,j,padding};
                        h1InSeedSet[161]<={hashValue[80][255:0],salt,t,j,padding};
                        h1InSeedSet[162]<={hashValue[81][511:256],salt,t,j,padding};
                        h1InSeedSet[163]<={hashValue[81][255:0],salt,t,j,padding};
                        h1InSeedSet[164]<={hashValue[82][511:256],salt,t,j,padding};
                        h1InSeedSet[165]<={hashValue[82][255:0],salt,t,j,padding};
                        h1InSeedSet[166]<={hashValue[83][511:256],salt,t,j,padding};
                        h1InSeedSet[167]<={hashValue[83][255:0],salt,t,j,padding};
                        h1InSeedSet[168]<={hashValue[84][511:256],salt,t,j,padding};
                        h1InSeedSet[169]<={hashValue[84][255:0],salt,t,j,padding};
                        h1InSeedSet[170]<={hashValue[85][511:256],salt,t,j,padding};
                        h1InSeedSet[171]<={hashValue[85][255:0],salt,t,j,padding};
                        h1InSeedSet[172]<={hashValue[86][511:256],salt,t,j,padding};
                        h1InSeedSet[173]<={hashValue[86][255:0],salt,t,j,padding};
                        h1InSeedSet[174]<={hashValue[87][511:256],salt,t,j,padding};
                        h1InSeedSet[175]<={hashValue[87][255:0],salt,t,j,padding};
                        h1InSeedSet[176]<={hashValue[88][511:256],salt,t,j,padding};
                        h1InSeedSet[177]<={hashValue[88][255:0],salt,t,j,padding};
                        h1InSeedSet[178]<={hashValue[89][511:256],salt,t,j,padding};
                        h1InSeedSet[179]<={hashValue[89][255:0],salt,t,j,padding};
                        h1InSeedSet[180]<={hashValue[90][511:256],salt,t,j,padding};
                        h1InSeedSet[181]<={hashValue[90][255:0],salt,t,j,padding};
                        h1InSeedSet[182]<={hashValue[91][511:256],salt,t,j,padding};
                        h1InSeedSet[183]<={hashValue[91][255:0],salt,t,j,padding};
                        h1InSeedSet[184]<={hashValue[92][511:256],salt,t,j,padding};
                        h1InSeedSet[185]<={hashValue[92][255:0],salt,t,j,padding};
                        h1InSeedSet[186]<={hashValue[93][511:256],salt,t,j,padding};
                        h1InSeedSet[187]<={hashValue[93][255:0],salt,t,j,padding};
                        h1InSeedSet[188]<={hashValue[94][511:256],salt,t,j,padding};
                        h1InSeedSet[189]<={hashValue[94][255:0],salt,t,j,padding};
                        h1InSeedSet[190]<={hashValue[95][511:256],salt,t,j,padding};
                        h1InSeedSet[191]<={hashValue[95][255:0],salt,t,j,padding};
                        h1InSeedSet[192]<={hashValue[96][511:256],salt,t,j,padding};
                        h1InSeedSet[193]<={hashValue[96][255:0],salt,t,j,padding};
                        h1InSeedSet[194]<={hashValue[97][511:256],salt,t,j,padding};
                        h1InSeedSet[195]<={hashValue[97][255:0],salt,t,j,padding};
                        h1InSeedSet[196]<={hashValue[98][511:256],salt,t,j,padding};
                        h1InSeedSet[197]<={hashValue[98][255:0],salt,t,j,padding};
                        h1InSeedSet[198]<={hashValue[99][511:256],salt,t,j,padding};
                        h1InSeedSet[199]<={hashValue[99][255:0],salt,t,j,padding};
                        h1InSeedSet[200]<={hashValue[100][511:256],salt,t,j,padding};
                        h1InSeedSet[201]<={hashValue[100][255:0],salt,t,j,padding};
                        h1InSeedSet[202]<={hashValue[101][511:256],salt,t,j,padding};
                        h1InSeedSet[203]<={hashValue[101][255:0],salt,t,j,padding};
                        h1InSeedSet[204]<={hashValue[102][511:256],salt,t,j,padding};
                        h1InSeedSet[205]<={hashValue[102][255:0],salt,t,j,padding};
                        h1InSeedSet[206]<={hashValue[103][511:256],salt,t,j,padding};
                        h1InSeedSet[207]<={hashValue[103][255:0],salt,t,j,padding};
                        h1InSeedSet[208]<={hashValue[104][511:256],salt,t,j,padding};
                        h1InSeedSet[209]<={hashValue[104][255:0],salt,t,j,padding};
                        h1InSeedSet[210]<={hashValue[105][511:256],salt,t,j,padding};
                        h1InSeedSet[211]<={hashValue[105][255:0],salt,t,j,padding};
                        h1InSeedSet[212]<={hashValue[106][511:256],salt,t,j,padding};
                        h1InSeedSet[213]<={hashValue[106][255:0],salt,t,j,padding};
                        h1InSeedSet[214]<={hashValue[107][511:256],salt,t,j,padding};
                        h1InSeedSet[215]<={hashValue[107][255:0],salt,t,j,padding};
                        h1InSeedSet[216]<={hashValue[108][511:256],salt,t,j,padding};
                        h1InSeedSet[217]<={hashValue[108][255:0],salt,t,j,padding};
                        h1InSeedSet[218]<={hashValue[109][511:256],salt,t,j,padding};
                        h1InSeedSet[219]<={hashValue[109][255:0],salt,t,j,padding};
                        h1InSeedSet[220]<={hashValue[110][511:256],salt,t,j,padding};
                        h1InSeedSet[221]<={hashValue[110][255:0],salt,t,j,padding};
                        h1InSeedSet[222]<={hashValue[111][511:256],salt,t,j,padding};
                        h1InSeedSet[223]<={hashValue[111][255:0],salt,t,j,padding};
                        h1InSeedSet[224]<={hashValue[112][511:256],salt,t,j,padding};
                        h1InSeedSet[225]<={hashValue[112][255:0],salt,t,j,padding};
                        h1InSeedSet[226]<={hashValue[113][511:256],salt,t,j,padding};
                        h1InSeedSet[227]<={hashValue[113][255:0],salt,t,j,padding};
                        h1InSeedSet[228]<={hashValue[114][511:256],salt,t,j,padding};
                        h1InSeedSet[229]<={hashValue[114][255:0],salt,t,j,padding};
                        h1InSeedSet[230]<={hashValue[115][511:256],salt,t,j,padding};
                        h1InSeedSet[231]<={hashValue[115][255:0],salt,t,j,padding};
                        h1InSeedSet[232]<={hashValue[116][511:256],salt,t,j,padding};
                        h1InSeedSet[233]<={hashValue[116][255:0],salt,t,j,padding};
                        h1InSeedSet[234]<={hashValue[117][511:256],salt,t,j,padding};
                        h1InSeedSet[235]<={hashValue[117][255:0],salt,t,j,padding};
                        h1InSeedSet[236]<={hashValue[118][511:256],salt,t,j,padding};
                        h1InSeedSet[237]<={hashValue[118][255:0],salt,t,j,padding};
                        h1InSeedSet[238]<={hashValue[119][511:256],salt,t,j,padding};
                        h1InSeedSet[239]<={hashValue[119][255:0],salt,t,j,padding};
                        h1InSeedSet[240]<={hashValue[120][511:256],salt,t,j,padding};
                        h1InSeedSet[241]<={hashValue[120][255:0],salt,t,j,padding};
                        h1InSeedSet[242]<={hashValue[121][511:256],salt,t,j,padding};
                        h1InSeedSet[243]<={hashValue[121][255:0],salt,t,j,padding};
                        h1InSeedSet[244]<={hashValue[122][511:256],salt,t,j,padding};
                        h1InSeedSet[245]<={hashValue[122][255:0],salt,t,j,padding};
                        h1InSeedSet[246]<={hashValue[123][511:256],salt,t,j,padding};
                        h1InSeedSet[247]<={hashValue[123][255:0],salt,t,j,padding};
                        h1InSeedSet[248]<={hashValue[124][511:256],salt,t,j,padding};
                        h1InSeedSet[249]<={hashValue[124][255:0],salt,t,j,padding};
                        h1InSeedSet[250]<={hashValue[125][511:256],salt,t,j,padding};
                        h1InSeedSet[251]<={hashValue[125][255:0],salt,t,j,padding};
                        h1InSeedSet[252]<={hashValue[126][511:256],salt,t,j,padding};
                        h1InSeedSet[253]<={hashValue[126][255:0],salt,t,j,padding};
                        h1InSeedSet[254]<={hashValue[127][511:256],salt,t,j,padding};
                        h1InSeedSet[255]<={hashValue[127][255:0],salt,t,j,padding};
                        h1InSeedSet[256]<={hashValue[128][511:256],salt,t,j,padding};
                        h1InSeedSet[257]<={hashValue[128][255:0],salt,t,j,padding};
                        h1InSeedSet[258]<={hashValue[129][511:256],salt,t,j,padding};
                        h1InSeedSet[259]<={hashValue[129][255:0],salt,t,j,padding};
                        h1InSeedSet[260]<={hashValue[130][511:256],salt,t,j,padding};
                        h1InSeedSet[261]<={hashValue[130][255:0],salt,t,j,padding};
                        h1InSeedSet[262]<={hashValue[131][511:256],salt,t,j,padding};
                        h1InSeedSet[263]<={hashValue[131][255:0],salt,t,j,padding};
                        h1InSeedSet[264]<={hashValue[132][511:256],salt,t,j,padding};
                        h1InSeedSet[265]<={hashValue[132][255:0],salt,t,j,padding};
                        h1InSeedSet[266]<={hashValue[133][511:256],salt,t,j,padding};
                        h1InSeedSet[267]<={hashValue[133][255:0],salt,t,j,padding};
                        h1InSeedSet[268]<={hashValue[134][511:256],salt,t,j,padding};
                        h1InSeedSet[269]<={hashValue[134][255:0],salt,t,j,padding};
                        h1InSeedSet[270]<={hashValue[135][511:256],salt,t,j,padding};
                        h1InSeedSet[271]<={hashValue[135][255:0],salt,t,j,padding};
                        h1InSeedSet[272]<={hashValue[136][511:256],salt,t,j,padding};
                        h1InSeedSet[273]<={hashValue[136][255:0],salt,t,j,padding};
                        h1InSeedSet[274]<={hashValue[137][511:256],salt,t,j,padding};
                        h1InSeedSet[275]<={hashValue[137][255:0],salt,t,j,padding};
                        h1InSeedSet[276]<={hashValue[138][511:256],salt,t,j,padding};
                        h1InSeedSet[277]<={hashValue[138][255:0],salt,t,j,padding};
                        h1InSeedSet[278]<={hashValue[139][511:256],salt,t,j,padding};
                        h1InSeedSet[279]<={hashValue[139][255:0],salt,t,j,padding};
                        h1InSeedSet[280]<={hashValue[140][511:256],salt,t,j,padding};
                        h1InSeedSet[281]<={hashValue[140][255:0],salt,t,j,padding};
                        h1InSeedSet[282]<={hashValue[141][511:256],salt,t,j,padding};
                        h1InSeedSet[283]<={hashValue[141][255:0],salt,t,j,padding};
                        h1InSeedSet[284]<={hashValue[142][511:256],salt,t,j,padding};
                        h1InSeedSet[285]<={hashValue[142][255:0],salt,t,j,padding};
                        h1InSeedSet[286]<={hashValue[143][511:256],salt,t,j,padding};
                        h1InSeedSet[287]<={hashValue[143][255:0],salt,t,j,padding};
                        h1InSeedSet[288]<={hashValue[144][511:256],salt,t,j,padding};
                        h1InSeedSet[289]<={hashValue[144][255:0],salt,t,j,padding};
                        h1InSeedSet[290]<={hashValue[145][511:256],salt,t,j,padding};
                        h1InSeedSet[291]<={hashValue[145][255:0],salt,t,j,padding};
                        h1InSeedSet[292]<={hashValue[146][511:256],salt,t,j,padding};
                        h1InSeedSet[293]<={hashValue[146][255:0],salt,t,j,padding};
                        h1InSeedSet[294]<={hashValue[147][511:256],salt,t,j,padding};
                        h1InSeedSet[295]<={hashValue[147][255:0],salt,t,j,padding};
                        h1InSeedSet[296]<={hashValue[148][511:256],salt,t,j,padding};
                        h1InSeedSet[297]<={hashValue[148][255:0],salt,t,j,padding};
                        h1InSeedSet[298]<={hashValue[149][511:256],salt,t,j,padding};
                        h1InSeedSet[299]<={hashValue[149][255:0],salt,t,j,padding};
                        h1InSeedSet[300]<={hashValue[150][511:256],salt,t,j,padding};
                        
                    end
                                   
            end
            if(state==2) begin
                iseed[154111:153600] <= hashValue[0];
                iseed[153599:153088] <= hashValue[1];
                iseed[153087:152576] <= hashValue[2];
                iseed[152575:152064] <= hashValue[3];
                iseed[152063:151552] <= hashValue[4];
                iseed[151551:151040] <= hashValue[5];
                iseed[151039:150528] <= hashValue[6];
                iseed[150527:150016] <= hashValue[7];
                iseed[150015:149504] <= hashValue[8];
                iseed[149503:148992] <= hashValue[9];
                iseed[148991:148480] <= hashValue[10];
                iseed[148479:147968] <= hashValue[11];
                iseed[147967:147456] <= hashValue[12];
                iseed[147455:146944] <= hashValue[13];
                iseed[146943:146432] <= hashValue[14];
                iseed[146431:145920] <= hashValue[15];
                iseed[145919:145408] <= hashValue[16];
                iseed[145407:144896] <= hashValue[17];
                iseed[144895:144384] <= hashValue[18];
                iseed[144383:143872] <= hashValue[19];
                iseed[143871:143360] <= hashValue[20];
                iseed[143359:142848] <= hashValue[21];
                iseed[142847:142336] <= hashValue[22];
                iseed[142335:141824] <= hashValue[23];
                iseed[141823:141312] <= hashValue[24];
                iseed[141311:140800] <= hashValue[25];
                iseed[140799:140288] <= hashValue[26];
                iseed[140287:139776] <= hashValue[27];
                iseed[139775:139264] <= hashValue[28];
                iseed[139263:138752] <= hashValue[29];
                iseed[138751:138240] <= hashValue[30];
                iseed[138239:137728] <= hashValue[31];
                iseed[137727:137216] <= hashValue[32];
                iseed[137215:136704] <= hashValue[33];
                iseed[136703:136192] <= hashValue[34];
                iseed[136191:135680] <= hashValue[35];
                iseed[135679:135168] <= hashValue[36];
                iseed[135167:134656] <= hashValue[37];
                iseed[134655:134144] <= hashValue[38];
                iseed[134143:133632] <= hashValue[39];
                iseed[133631:133120] <= hashValue[40];
                iseed[133119:132608] <= hashValue[41];
                iseed[132607:132096] <= hashValue[42];
                iseed[132095:131584] <= hashValue[43];
                iseed[131583:131072] <= hashValue[44];
                iseed[131071:130560] <= hashValue[45];
                iseed[130559:130048] <= hashValue[46];
                iseed[130047:129536] <= hashValue[47];
                iseed[129535:129024] <= hashValue[48];
                iseed[129023:128512] <= hashValue[49];
                iseed[128511:128000] <= hashValue[50];
                iseed[127999:127488] <= hashValue[51];
                iseed[127487:126976] <= hashValue[52];
                iseed[126975:126464] <= hashValue[53];
                iseed[126463:125952] <= hashValue[54];
                iseed[125951:125440] <= hashValue[55];
                iseed[125439:124928] <= hashValue[56];
                iseed[124927:124416] <= hashValue[57];
                iseed[124415:123904] <= hashValue[58];
                iseed[123903:123392] <= hashValue[59];
                iseed[123391:122880] <= hashValue[60];
                iseed[122879:122368] <= hashValue[61];
                iseed[122367:121856] <= hashValue[62];
                iseed[121855:121344] <= hashValue[63];
                iseed[121343:120832] <= hashValue[64];
                iseed[120831:120320] <= hashValue[65];
                iseed[120319:119808] <= hashValue[66];
                iseed[119807:119296] <= hashValue[67];
                iseed[119295:118784] <= hashValue[68];
                iseed[118783:118272] <= hashValue[69];
                iseed[118271:117760] <= hashValue[70];
                iseed[117759:117248] <= hashValue[71];
                iseed[117247:116736] <= hashValue[72];
                iseed[116735:116224] <= hashValue[73];
                iseed[116223:115712] <= hashValue[74];
                iseed[115711:115200] <= hashValue[75];
                iseed[115199:114688] <= hashValue[76];
                iseed[114687:114176] <= hashValue[77];
                iseed[114175:113664] <= hashValue[78];
                iseed[113663:113152] <= hashValue[79];
                iseed[113151:112640] <= hashValue[80];
                iseed[112639:112128] <= hashValue[81];
                iseed[112127:111616] <= hashValue[82];
                iseed[111615:111104] <= hashValue[83];
                iseed[111103:110592] <= hashValue[84];
                iseed[110591:110080] <= hashValue[85];
                iseed[110079:109568] <= hashValue[86];
                iseed[109567:109056] <= hashValue[87];
                iseed[109055:108544] <= hashValue[88];
                iseed[108543:108032] <= hashValue[89];
                iseed[108031:107520] <= hashValue[90];
                iseed[107519:107008] <= hashValue[91];
                iseed[107007:106496] <= hashValue[92];
                iseed[106495:105984] <= hashValue[93];
                iseed[105983:105472] <= hashValue[94];
                iseed[105471:104960] <= hashValue[95];
                iseed[104959:104448] <= hashValue[96];
                iseed[104447:103936] <= hashValue[97];
                iseed[103935:103424] <= hashValue[98];
                iseed[103423:102912] <= hashValue[99];
                iseed[102911:102400] <= hashValue[100];
                iseed[102399:101888] <= hashValue[101];
                iseed[101887:101376] <= hashValue[102];
                iseed[101375:100864] <= hashValue[103];
                iseed[100863:100352] <= hashValue[104];
                iseed[100351:99840] <= hashValue[105];
                iseed[99839:99328] <= hashValue[106];
                iseed[99327:98816] <= hashValue[107];
                iseed[98815:98304] <= hashValue[108];
                iseed[98303:97792] <= hashValue[109];
                iseed[97791:97280] <= hashValue[110];
                iseed[97279:96768] <= hashValue[111];
                iseed[96767:96256] <= hashValue[112];
                iseed[96255:95744] <= hashValue[113];
                iseed[95743:95232] <= hashValue[114];
                iseed[95231:94720] <= hashValue[115];
                iseed[94719:94208] <= hashValue[116];
                iseed[94207:93696] <= hashValue[117];
                iseed[93695:93184] <= hashValue[118];
                iseed[93183:92672] <= hashValue[119];
                iseed[92671:92160] <= hashValue[120];
                iseed[92159:91648] <= hashValue[121];
                iseed[91647:91136] <= hashValue[122];
                iseed[91135:90624] <= hashValue[123];
                iseed[90623:90112] <= hashValue[124];
                iseed[90111:89600] <= hashValue[125];
                iseed[89599:89088] <= hashValue[126];
                iseed[89087:88576] <= hashValue[127];
                iseed[88575:88064] <= hashValue[128];
                iseed[88063:87552] <= hashValue[129];
                iseed[87551:87040] <= hashValue[130];
                iseed[87039:86528] <= hashValue[131];
                iseed[86527:86016] <= hashValue[132];
                iseed[86015:85504] <= hashValue[133];
                iseed[85503:84992] <= hashValue[134];
                iseed[84991:84480] <= hashValue[135];
                iseed[84479:83968] <= hashValue[136];
                iseed[83967:83456] <= hashValue[137];
                iseed[83455:82944] <= hashValue[138];
                iseed[82943:82432] <= hashValue[139];
                iseed[82431:81920] <= hashValue[140];
                iseed[81919:81408] <= hashValue[141];
                iseed[81407:80896] <= hashValue[142];
                iseed[80895:80384] <= hashValue[143];
                iseed[80383:79872] <= hashValue[144];
                iseed[79871:79360] <= hashValue[145];
                iseed[79359:78848] <= hashValue[146];
                iseed[78847:78336] <= hashValue[147];
                iseed[78335:77824] <= hashValue[148];
                iseed[77823:77312] <= hashValue[149];
                iseed[77311:76800] <= hashValue[150];
                iseed[76799:76288] <= hashValue[151];
                iseed[76287:75776] <= hashValue[152];
                iseed[75775:75264] <= hashValue[153];
                iseed[75263:74752] <= hashValue[154];
                iseed[74751:74240] <= hashValue[155];
                iseed[74239:73728] <= hashValue[156];
                iseed[73727:73216] <= hashValue[157];
                iseed[73215:72704] <= hashValue[158];
                iseed[72703:72192] <= hashValue[159];
                iseed[72191:71680] <= hashValue[160];
                iseed[71679:71168] <= hashValue[161];
                iseed[71167:70656] <= hashValue[162];
                iseed[70655:70144] <= hashValue[163];
                iseed[70143:69632] <= hashValue[164];
                iseed[69631:69120] <= hashValue[165];
                iseed[69119:68608] <= hashValue[166];
                iseed[68607:68096] <= hashValue[167];
                iseed[68095:67584] <= hashValue[168];
                iseed[67583:67072] <= hashValue[169];
                iseed[67071:66560] <= hashValue[170];
                iseed[66559:66048] <= hashValue[171];
                iseed[66047:65536] <= hashValue[172];
                iseed[65535:65024] <= hashValue[173];
                iseed[65023:64512] <= hashValue[174];
                iseed[64511:64000] <= hashValue[175];
                iseed[63999:63488] <= hashValue[176];
                iseed[63487:62976] <= hashValue[177];
                iseed[62975:62464] <= hashValue[178];
                iseed[62463:61952] <= hashValue[179];
                iseed[61951:61440] <= hashValue[180];
                iseed[61439:60928] <= hashValue[181];
                iseed[60927:60416] <= hashValue[182];
                iseed[60415:59904] <= hashValue[183];
                iseed[59903:59392] <= hashValue[184];
                iseed[59391:58880] <= hashValue[185];
                iseed[58879:58368] <= hashValue[186];
                iseed[58367:57856] <= hashValue[187];
                iseed[57855:57344] <= hashValue[188];
                iseed[57343:56832] <= hashValue[189];
                iseed[56831:56320] <= hashValue[190];
                iseed[56319:55808] <= hashValue[191];
                iseed[55807:55296] <= hashValue[192];
                iseed[55295:54784] <= hashValue[193];
                iseed[54783:54272] <= hashValue[194];
                iseed[54271:53760] <= hashValue[195];
                iseed[53759:53248] <= hashValue[196];
                iseed[53247:52736] <= hashValue[197];
                iseed[52735:52224] <= hashValue[198];
                iseed[52223:51712] <= hashValue[199];
                iseed[51711:51200] <= hashValue[200];
                iseed[51199:50688] <= hashValue[201];
                iseed[50687:50176] <= hashValue[202];
                iseed[50175:49664] <= hashValue[203];
                iseed[49663:49152] <= hashValue[204];
                iseed[49151:48640] <= hashValue[205];
                iseed[48639:48128] <= hashValue[206];
                iseed[48127:47616] <= hashValue[207];
                iseed[47615:47104] <= hashValue[208];
                iseed[47103:46592] <= hashValue[209];
                iseed[46591:46080] <= hashValue[210];
                iseed[46079:45568] <= hashValue[211];
                iseed[45567:45056] <= hashValue[212];
                iseed[45055:44544] <= hashValue[213];
                iseed[44543:44032] <= hashValue[214];
                iseed[44031:43520] <= hashValue[215];
                iseed[43519:43008] <= hashValue[216];
                iseed[43007:42496] <= hashValue[217];
                iseed[42495:41984] <= hashValue[218];
                iseed[41983:41472] <= hashValue[219];
                iseed[41471:40960] <= hashValue[220];
                iseed[40959:40448] <= hashValue[221];
                iseed[40447:39936] <= hashValue[222];
                iseed[39935:39424] <= hashValue[223];
                iseed[39423:38912] <= hashValue[224];
                iseed[38911:38400] <= hashValue[225];
                iseed[38399:37888] <= hashValue[226];
                iseed[37887:37376] <= hashValue[227];
                iseed[37375:36864] <= hashValue[228];
                iseed[36863:36352] <= hashValue[229];
                iseed[36351:35840] <= hashValue[230];
                iseed[35839:35328] <= hashValue[231];
                iseed[35327:34816] <= hashValue[232];
                iseed[34815:34304] <= hashValue[233];
                iseed[34303:33792] <= hashValue[234];
                iseed[33791:33280] <= hashValue[235];
                iseed[33279:32768] <= hashValue[236];
                iseed[32767:32256] <= hashValue[237];
                iseed[32255:31744] <= hashValue[238];
                iseed[31743:31232] <= hashValue[239];
                iseed[31231:30720] <= hashValue[240];
                iseed[30719:30208] <= hashValue[241];
                iseed[30207:29696] <= hashValue[242];
                iseed[29695:29184] <= hashValue[243];
                iseed[29183:28672] <= hashValue[244];
                iseed[28671:28160] <= hashValue[245];
                iseed[28159:27648] <= hashValue[246];
                iseed[27647:27136] <= hashValue[247];
                iseed[27135:26624] <= hashValue[248];
                iseed[26623:26112] <= hashValue[249];
                iseed[26111:25600] <= hashValue[250];
                iseed[25599:25088] <= hashValue[251];
                iseed[25087:24576] <= hashValue[252];
                iseed[24575:24064] <= hashValue[253];
                iseed[24063:23552] <= hashValue[254];
                iseed[23551:23040] <= hashValue[255];
                iseed[23039:22528] <= hashValue[256];
                iseed[22527:22016] <= hashValue[257];
                iseed[22015:21504] <= hashValue[258];
                iseed[21503:20992] <= hashValue[259];
                iseed[20991:20480] <= hashValue[260];
                iseed[20479:19968] <= hashValue[261];
                iseed[19967:19456] <= hashValue[262];
                iseed[19455:18944] <= hashValue[263];
                iseed[18943:18432] <= hashValue[264];
                iseed[18431:17920] <= hashValue[265];
                iseed[17919:17408] <= hashValue[266];
                iseed[17407:16896] <= hashValue[267];
                iseed[16895:16384] <= hashValue[268];
                iseed[16383:15872] <= hashValue[269];
                iseed[15871:15360] <= hashValue[270];
                iseed[15359:14848] <= hashValue[271];
                iseed[14847:14336] <= hashValue[272];
                iseed[14335:13824] <= hashValue[273];
                iseed[13823:13312] <= hashValue[274];
                iseed[13311:12800] <= hashValue[275];
                iseed[12799:12288] <= hashValue[276];
                iseed[12287:11776] <= hashValue[277];
                iseed[11775:11264] <= hashValue[278];
                iseed[11263:10752] <= hashValue[279];
                iseed[10751:10240] <= hashValue[280];
                iseed[10239:9728] <= hashValue[281];
                iseed[9727:9216] <= hashValue[282];
                iseed[9215:8704] <= hashValue[283];
                iseed[8703:8192] <= hashValue[284];
                iseed[8191:7680] <= hashValue[285];
                iseed[7679:7168] <= hashValue[286];
                iseed[7167:6656] <= hashValue[287];
                iseed[6655:6144] <= hashValue[288];
                iseed[6143:5632] <= hashValue[289];
                iseed[5631:5120] <= hashValue[290];
                iseed[5119:4608] <= hashValue[291];
                iseed[4607:4096] <= hashValue[292];
                iseed[4095:3584] <= hashValue[293];
                iseed[3583:3072] <= hashValue[294];
                iseed[3071:2560] <= hashValue[295];
                iseed[2559:2048] <= hashValue[296];
                iseed[2047:1536] <= hashValue[297];
                iseed[1535:1024] <= hashValue[298];
                iseed[1023:512] <= hashValue[299];
                iseed[511:0] <= hashValue[300];
                tree_set_end<=1;
                state <= 3;
            end
            if(state==3) begin
                tree_set_end <= 0;
                state<=0;
            end
        end

    end

    

H h0(clk,reset,0,h1InSeedSet[0],0,Hstart[0],restart[0],groupNum,hashValue[0],en_end[0]);
H h1(clk,reset,0,h1InSeedSet[1],0,Hstart[1],restart[1],groupNum,hashValue[1],en_end[1]);
H h2(clk,reset,0,h1InSeedSet[2],0,Hstart[2],restart[2],groupNum,hashValue[2],en_end[2]);
H h3(clk,reset,0,h1InSeedSet[3],0,Hstart[3],restart[3],groupNum,hashValue[3],en_end[3]);
H h4(clk,reset,0,h1InSeedSet[4],0,Hstart[4],restart[4],groupNum,hashValue[4],en_end[4]);
H h5(clk,reset,0,h1InSeedSet[5],0,Hstart[5],restart[5],groupNum,hashValue[5],en_end[5]);
H h6(clk,reset,0,h1InSeedSet[6],0,Hstart[6],restart[6],groupNum,hashValue[6],en_end[6]);
H h7(clk,reset,0,h1InSeedSet[7],0,Hstart[7],restart[7],groupNum,hashValue[7],en_end[7]);
H h8(clk,reset,0,h1InSeedSet[8],0,Hstart[8],restart[8],groupNum,hashValue[8],en_end[8]);
H h9(clk,reset,0,h1InSeedSet[9],0,Hstart[9],restart[9],groupNum,hashValue[9],en_end[9]);
H h10(clk,reset,0,h1InSeedSet[10],0,Hstart[10],restart[10],groupNum,hashValue[10],en_end[10]);
H h11(clk,reset,0,h1InSeedSet[11],0,Hstart[11],restart[11],groupNum,hashValue[11],en_end[11]);
H h12(clk,reset,0,h1InSeedSet[12],0,Hstart[12],restart[12],groupNum,hashValue[12],en_end[12]);
H h13(clk,reset,0,h1InSeedSet[13],0,Hstart[13],restart[13],groupNum,hashValue[13],en_end[13]);
H h14(clk,reset,0,h1InSeedSet[14],0,Hstart[14],restart[14],groupNum,hashValue[14],en_end[14]);
H h15(clk,reset,0,h1InSeedSet[15],0,Hstart[15],restart[15],groupNum,hashValue[15],en_end[15]);
H h16(clk,reset,0,h1InSeedSet[16],0,Hstart[16],restart[16],groupNum,hashValue[16],en_end[16]);
H h17(clk,reset,0,h1InSeedSet[17],0,Hstart[17],restart[17],groupNum,hashValue[17],en_end[17]);
H h18(clk,reset,0,h1InSeedSet[18],0,Hstart[18],restart[18],groupNum,hashValue[18],en_end[18]);
H h19(clk,reset,0,h1InSeedSet[19],0,Hstart[19],restart[19],groupNum,hashValue[19],en_end[19]);
H h20(clk,reset,0,h1InSeedSet[20],0,Hstart[20],restart[20],groupNum,hashValue[20],en_end[20]);
H h21(clk,reset,0,h1InSeedSet[21],0,Hstart[21],restart[21],groupNum,hashValue[21],en_end[21]);
H h22(clk,reset,0,h1InSeedSet[22],0,Hstart[22],restart[22],groupNum,hashValue[22],en_end[22]);
H h23(clk,reset,0,h1InSeedSet[23],0,Hstart[23],restart[23],groupNum,hashValue[23],en_end[23]);
H h24(clk,reset,0,h1InSeedSet[24],0,Hstart[24],restart[24],groupNum,hashValue[24],en_end[24]);
H h25(clk,reset,0,h1InSeedSet[25],0,Hstart[25],restart[25],groupNum,hashValue[25],en_end[25]);
H h26(clk,reset,0,h1InSeedSet[26],0,Hstart[26],restart[26],groupNum,hashValue[26],en_end[26]);
H h27(clk,reset,0,h1InSeedSet[27],0,Hstart[27],restart[27],groupNum,hashValue[27],en_end[27]);
H h28(clk,reset,0,h1InSeedSet[28],0,Hstart[28],restart[28],groupNum,hashValue[28],en_end[28]);
H h29(clk,reset,0,h1InSeedSet[29],0,Hstart[29],restart[29],groupNum,hashValue[29],en_end[29]);
H h30(clk,reset,0,h1InSeedSet[30],0,Hstart[30],restart[30],groupNum,hashValue[30],en_end[30]);
H h31(clk,reset,0,h1InSeedSet[31],0,Hstart[31],restart[31],groupNum,hashValue[31],en_end[31]);
H h32(clk,reset,0,h1InSeedSet[32],0,Hstart[32],restart[32],groupNum,hashValue[32],en_end[32]);
H h33(clk,reset,0,h1InSeedSet[33],0,Hstart[33],restart[33],groupNum,hashValue[33],en_end[33]);
H h34(clk,reset,0,h1InSeedSet[34],0,Hstart[34],restart[34],groupNum,hashValue[34],en_end[34]);
H h35(clk,reset,0,h1InSeedSet[35],0,Hstart[35],restart[35],groupNum,hashValue[35],en_end[35]);
H h36(clk,reset,0,h1InSeedSet[36],0,Hstart[36],restart[36],groupNum,hashValue[36],en_end[36]);
H h37(clk,reset,0,h1InSeedSet[37],0,Hstart[37],restart[37],groupNum,hashValue[37],en_end[37]);
H h38(clk,reset,0,h1InSeedSet[38],0,Hstart[38],restart[38],groupNum,hashValue[38],en_end[38]);
H h39(clk,reset,0,h1InSeedSet[39],0,Hstart[39],restart[39],groupNum,hashValue[39],en_end[39]);
H h40(clk,reset,0,h1InSeedSet[40],0,Hstart[40],restart[40],groupNum,hashValue[40],en_end[40]);
H h41(clk,reset,0,h1InSeedSet[41],0,Hstart[41],restart[41],groupNum,hashValue[41],en_end[41]);
H h42(clk,reset,0,h1InSeedSet[42],0,Hstart[42],restart[42],groupNum,hashValue[42],en_end[42]);
H h43(clk,reset,0,h1InSeedSet[43],0,Hstart[43],restart[43],groupNum,hashValue[43],en_end[43]);
H h44(clk,reset,0,h1InSeedSet[44],0,Hstart[44],restart[44],groupNum,hashValue[44],en_end[44]);
H h45(clk,reset,0,h1InSeedSet[45],0,Hstart[45],restart[45],groupNum,hashValue[45],en_end[45]);
H h46(clk,reset,0,h1InSeedSet[46],0,Hstart[46],restart[46],groupNum,hashValue[46],en_end[46]);
H h47(clk,reset,0,h1InSeedSet[47],0,Hstart[47],restart[47],groupNum,hashValue[47],en_end[47]);
H h48(clk,reset,0,h1InSeedSet[48],0,Hstart[48],restart[48],groupNum,hashValue[48],en_end[48]);
H h49(clk,reset,0,h1InSeedSet[49],0,Hstart[49],restart[49],groupNum,hashValue[49],en_end[49]);
H h50(clk,reset,0,h1InSeedSet[50],0,Hstart[50],restart[50],groupNum,hashValue[50],en_end[50]);
H h51(clk,reset,0,h1InSeedSet[51],0,Hstart[51],restart[51],groupNum,hashValue[51],en_end[51]);
H h52(clk,reset,0,h1InSeedSet[52],0,Hstart[52],restart[52],groupNum,hashValue[52],en_end[52]);
H h53(clk,reset,0,h1InSeedSet[53],0,Hstart[53],restart[53],groupNum,hashValue[53],en_end[53]);
H h54(clk,reset,0,h1InSeedSet[54],0,Hstart[54],restart[54],groupNum,hashValue[54],en_end[54]);
H h55(clk,reset,0,h1InSeedSet[55],0,Hstart[55],restart[55],groupNum,hashValue[55],en_end[55]);
H h56(clk,reset,0,h1InSeedSet[56],0,Hstart[56],restart[56],groupNum,hashValue[56],en_end[56]);
H h57(clk,reset,0,h1InSeedSet[57],0,Hstart[57],restart[57],groupNum,hashValue[57],en_end[57]);
H h58(clk,reset,0,h1InSeedSet[58],0,Hstart[58],restart[58],groupNum,hashValue[58],en_end[58]);
H h59(clk,reset,0,h1InSeedSet[59],0,Hstart[59],restart[59],groupNum,hashValue[59],en_end[59]);
H h60(clk,reset,0,h1InSeedSet[60],0,Hstart[60],restart[60],groupNum,hashValue[60],en_end[60]);
H h61(clk,reset,0,h1InSeedSet[61],0,Hstart[61],restart[61],groupNum,hashValue[61],en_end[61]);
H h62(clk,reset,0,h1InSeedSet[62],0,Hstart[62],restart[62],groupNum,hashValue[62],en_end[62]);
H h63(clk,reset,0,h1InSeedSet[63],0,Hstart[63],restart[63],groupNum,hashValue[63],en_end[63]);
H h64(clk,reset,0,h1InSeedSet[64],0,Hstart[64],restart[64],groupNum,hashValue[64],en_end[64]);
H h65(clk,reset,0,h1InSeedSet[65],0,Hstart[65],restart[65],groupNum,hashValue[65],en_end[65]);
H h66(clk,reset,0,h1InSeedSet[66],0,Hstart[66],restart[66],groupNum,hashValue[66],en_end[66]);
H h67(clk,reset,0,h1InSeedSet[67],0,Hstart[67],restart[67],groupNum,hashValue[67],en_end[67]);
H h68(clk,reset,0,h1InSeedSet[68],0,Hstart[68],restart[68],groupNum,hashValue[68],en_end[68]);
H h69(clk,reset,0,h1InSeedSet[69],0,Hstart[69],restart[69],groupNum,hashValue[69],en_end[69]);
H h70(clk,reset,0,h1InSeedSet[70],0,Hstart[70],restart[70],groupNum,hashValue[70],en_end[70]);
H h71(clk,reset,0,h1InSeedSet[71],0,Hstart[71],restart[71],groupNum,hashValue[71],en_end[71]);
H h72(clk,reset,0,h1InSeedSet[72],0,Hstart[72],restart[72],groupNum,hashValue[72],en_end[72]);
H h73(clk,reset,0,h1InSeedSet[73],0,Hstart[73],restart[73],groupNum,hashValue[73],en_end[73]);
H h74(clk,reset,0,h1InSeedSet[74],0,Hstart[74],restart[74],groupNum,hashValue[74],en_end[74]);
H h75(clk,reset,0,h1InSeedSet[75],0,Hstart[75],restart[75],groupNum,hashValue[75],en_end[75]);
H h76(clk,reset,0,h1InSeedSet[76],0,Hstart[76],restart[76],groupNum,hashValue[76],en_end[76]);
H h77(clk,reset,0,h1InSeedSet[77],0,Hstart[77],restart[77],groupNum,hashValue[77],en_end[77]);
H h78(clk,reset,0,h1InSeedSet[78],0,Hstart[78],restart[78],groupNum,hashValue[78],en_end[78]);
H h79(clk,reset,0,h1InSeedSet[79],0,Hstart[79],restart[79],groupNum,hashValue[79],en_end[79]);
H h80(clk,reset,0,h1InSeedSet[80],0,Hstart[80],restart[80],groupNum,hashValue[80],en_end[80]);
H h81(clk,reset,0,h1InSeedSet[81],0,Hstart[81],restart[81],groupNum,hashValue[81],en_end[81]);
H h82(clk,reset,0,h1InSeedSet[82],0,Hstart[82],restart[82],groupNum,hashValue[82],en_end[82]);
H h83(clk,reset,0,h1InSeedSet[83],0,Hstart[83],restart[83],groupNum,hashValue[83],en_end[83]);
H h84(clk,reset,0,h1InSeedSet[84],0,Hstart[84],restart[84],groupNum,hashValue[84],en_end[84]);
H h85(clk,reset,0,h1InSeedSet[85],0,Hstart[85],restart[85],groupNum,hashValue[85],en_end[85]);
H h86(clk,reset,0,h1InSeedSet[86],0,Hstart[86],restart[86],groupNum,hashValue[86],en_end[86]);
H h87(clk,reset,0,h1InSeedSet[87],0,Hstart[87],restart[87],groupNum,hashValue[87],en_end[87]);
H h88(clk,reset,0,h1InSeedSet[88],0,Hstart[88],restart[88],groupNum,hashValue[88],en_end[88]);
H h89(clk,reset,0,h1InSeedSet[89],0,Hstart[89],restart[89],groupNum,hashValue[89],en_end[89]);
H h90(clk,reset,0,h1InSeedSet[90],0,Hstart[90],restart[90],groupNum,hashValue[90],en_end[90]);
H h91(clk,reset,0,h1InSeedSet[91],0,Hstart[91],restart[91],groupNum,hashValue[91],en_end[91]);
H h92(clk,reset,0,h1InSeedSet[92],0,Hstart[92],restart[92],groupNum,hashValue[92],en_end[92]);
H h93(clk,reset,0,h1InSeedSet[93],0,Hstart[93],restart[93],groupNum,hashValue[93],en_end[93]);
H h94(clk,reset,0,h1InSeedSet[94],0,Hstart[94],restart[94],groupNum,hashValue[94],en_end[94]);
H h95(clk,reset,0,h1InSeedSet[95],0,Hstart[95],restart[95],groupNum,hashValue[95],en_end[95]);
H h96(clk,reset,0,h1InSeedSet[96],0,Hstart[96],restart[96],groupNum,hashValue[96],en_end[96]);
H h97(clk,reset,0,h1InSeedSet[97],0,Hstart[97],restart[97],groupNum,hashValue[97],en_end[97]);
H h98(clk,reset,0,h1InSeedSet[98],0,Hstart[98],restart[98],groupNum,hashValue[98],en_end[98]);
H h99(clk,reset,0,h1InSeedSet[99],0,Hstart[99],restart[99],groupNum,hashValue[99],en_end[99]);
H h100(clk,reset,0,h1InSeedSet[100],0,Hstart[100],restart[100],groupNum,hashValue[100],en_end[100]);
H h101(clk,reset,0,h1InSeedSet[101],0,Hstart[101],restart[101],groupNum,hashValue[101],en_end[101]);
H h102(clk,reset,0,h1InSeedSet[102],0,Hstart[102],restart[102],groupNum,hashValue[102],en_end[102]);
H h103(clk,reset,0,h1InSeedSet[103],0,Hstart[103],restart[103],groupNum,hashValue[103],en_end[103]);
H h104(clk,reset,0,h1InSeedSet[104],0,Hstart[104],restart[104],groupNum,hashValue[104],en_end[104]);
H h105(clk,reset,0,h1InSeedSet[105],0,Hstart[105],restart[105],groupNum,hashValue[105],en_end[105]);
H h106(clk,reset,0,h1InSeedSet[106],0,Hstart[106],restart[106],groupNum,hashValue[106],en_end[106]);
H h107(clk,reset,0,h1InSeedSet[107],0,Hstart[107],restart[107],groupNum,hashValue[107],en_end[107]);
H h108(clk,reset,0,h1InSeedSet[108],0,Hstart[108],restart[108],groupNum,hashValue[108],en_end[108]);
H h109(clk,reset,0,h1InSeedSet[109],0,Hstart[109],restart[109],groupNum,hashValue[109],en_end[109]);
H h110(clk,reset,0,h1InSeedSet[110],0,Hstart[110],restart[110],groupNum,hashValue[110],en_end[110]);
H h111(clk,reset,0,h1InSeedSet[111],0,Hstart[111],restart[111],groupNum,hashValue[111],en_end[111]);
H h112(clk,reset,0,h1InSeedSet[112],0,Hstart[112],restart[112],groupNum,hashValue[112],en_end[112]);
H h113(clk,reset,0,h1InSeedSet[113],0,Hstart[113],restart[113],groupNum,hashValue[113],en_end[113]);
H h114(clk,reset,0,h1InSeedSet[114],0,Hstart[114],restart[114],groupNum,hashValue[114],en_end[114]);
H h115(clk,reset,0,h1InSeedSet[115],0,Hstart[115],restart[115],groupNum,hashValue[115],en_end[115]);
H h116(clk,reset,0,h1InSeedSet[116],0,Hstart[116],restart[116],groupNum,hashValue[116],en_end[116]);
H h117(clk,reset,0,h1InSeedSet[117],0,Hstart[117],restart[117],groupNum,hashValue[117],en_end[117]);
H h118(clk,reset,0,h1InSeedSet[118],0,Hstart[118],restart[118],groupNum,hashValue[118],en_end[118]);
H h119(clk,reset,0,h1InSeedSet[119],0,Hstart[119],restart[119],groupNum,hashValue[119],en_end[119]);
H h120(clk,reset,0,h1InSeedSet[120],0,Hstart[120],restart[120],groupNum,hashValue[120],en_end[120]);
H h121(clk,reset,0,h1InSeedSet[121],0,Hstart[121],restart[121],groupNum,hashValue[121],en_end[121]);
H h122(clk,reset,0,h1InSeedSet[122],0,Hstart[122],restart[122],groupNum,hashValue[122],en_end[122]);
H h123(clk,reset,0,h1InSeedSet[123],0,Hstart[123],restart[123],groupNum,hashValue[123],en_end[123]);
H h124(clk,reset,0,h1InSeedSet[124],0,Hstart[124],restart[124],groupNum,hashValue[124],en_end[124]);
H h125(clk,reset,0,h1InSeedSet[125],0,Hstart[125],restart[125],groupNum,hashValue[125],en_end[125]);
H h126(clk,reset,0,h1InSeedSet[126],0,Hstart[126],restart[126],groupNum,hashValue[126],en_end[126]);
H h127(clk,reset,0,h1InSeedSet[127],0,Hstart[127],restart[127],groupNum,hashValue[127],en_end[127]);
H h128(clk,reset,0,h1InSeedSet[128],0,Hstart[128],restart[128],groupNum,hashValue[128],en_end[128]);
H h129(clk,reset,0,h1InSeedSet[129],0,Hstart[129],restart[129],groupNum,hashValue[129],en_end[129]);
H h130(clk,reset,0,h1InSeedSet[130],0,Hstart[130],restart[130],groupNum,hashValue[130],en_end[130]);
H h131(clk,reset,0,h1InSeedSet[131],0,Hstart[131],restart[131],groupNum,hashValue[131],en_end[131]);
H h132(clk,reset,0,h1InSeedSet[132],0,Hstart[132],restart[132],groupNum,hashValue[132],en_end[132]);
H h133(clk,reset,0,h1InSeedSet[133],0,Hstart[133],restart[133],groupNum,hashValue[133],en_end[133]);
H h134(clk,reset,0,h1InSeedSet[134],0,Hstart[134],restart[134],groupNum,hashValue[134],en_end[134]);
H h135(clk,reset,0,h1InSeedSet[135],0,Hstart[135],restart[135],groupNum,hashValue[135],en_end[135]);
H h136(clk,reset,0,h1InSeedSet[136],0,Hstart[136],restart[136],groupNum,hashValue[136],en_end[136]);
H h137(clk,reset,0,h1InSeedSet[137],0,Hstart[137],restart[137],groupNum,hashValue[137],en_end[137]);
H h138(clk,reset,0,h1InSeedSet[138],0,Hstart[138],restart[138],groupNum,hashValue[138],en_end[138]);
H h139(clk,reset,0,h1InSeedSet[139],0,Hstart[139],restart[139],groupNum,hashValue[139],en_end[139]);
H h140(clk,reset,0,h1InSeedSet[140],0,Hstart[140],restart[140],groupNum,hashValue[140],en_end[140]);
H h141(clk,reset,0,h1InSeedSet[141],0,Hstart[141],restart[141],groupNum,hashValue[141],en_end[141]);
H h142(clk,reset,0,h1InSeedSet[142],0,Hstart[142],restart[142],groupNum,hashValue[142],en_end[142]);
H h143(clk,reset,0,h1InSeedSet[143],0,Hstart[143],restart[143],groupNum,hashValue[143],en_end[143]);
H h144(clk,reset,0,h1InSeedSet[144],0,Hstart[144],restart[144],groupNum,hashValue[144],en_end[144]);
H h145(clk,reset,0,h1InSeedSet[145],0,Hstart[145],restart[145],groupNum,hashValue[145],en_end[145]);
H h146(clk,reset,0,h1InSeedSet[146],0,Hstart[146],restart[146],groupNum,hashValue[146],en_end[146]);
H h147(clk,reset,0,h1InSeedSet[147],0,Hstart[147],restart[147],groupNum,hashValue[147],en_end[147]);
H h148(clk,reset,0,h1InSeedSet[148],0,Hstart[148],restart[148],groupNum,hashValue[148],en_end[148]);
H h149(clk,reset,0,h1InSeedSet[149],0,Hstart[149],restart[149],groupNum,hashValue[149],en_end[149]);
H h150(clk,reset,0,h1InSeedSet[150],0,Hstart[150],restart[150],groupNum,hashValue[150],en_end[150]);
H h151(clk,reset,0,h1InSeedSet[151],0,Hstart[151],restart[151],groupNum,hashValue[151],en_end[151]);
H h152(clk,reset,0,h1InSeedSet[152],0,Hstart[152],restart[152],groupNum,hashValue[152],en_end[152]);
H h153(clk,reset,0,h1InSeedSet[153],0,Hstart[153],restart[153],groupNum,hashValue[153],en_end[153]);
H h154(clk,reset,0,h1InSeedSet[154],0,Hstart[154],restart[154],groupNum,hashValue[154],en_end[154]);
H h155(clk,reset,0,h1InSeedSet[155],0,Hstart[155],restart[155],groupNum,hashValue[155],en_end[155]);
H h156(clk,reset,0,h1InSeedSet[156],0,Hstart[156],restart[156],groupNum,hashValue[156],en_end[156]);
H h157(clk,reset,0,h1InSeedSet[157],0,Hstart[157],restart[157],groupNum,hashValue[157],en_end[157]);
H h158(clk,reset,0,h1InSeedSet[158],0,Hstart[158],restart[158],groupNum,hashValue[158],en_end[158]);
H h159(clk,reset,0,h1InSeedSet[159],0,Hstart[159],restart[159],groupNum,hashValue[159],en_end[159]);
H h160(clk,reset,0,h1InSeedSet[160],0,Hstart[160],restart[160],groupNum,hashValue[160],en_end[160]);
H h161(clk,reset,0,h1InSeedSet[161],0,Hstart[161],restart[161],groupNum,hashValue[161],en_end[161]);
H h162(clk,reset,0,h1InSeedSet[162],0,Hstart[162],restart[162],groupNum,hashValue[162],en_end[162]);
H h163(clk,reset,0,h1InSeedSet[163],0,Hstart[163],restart[163],groupNum,hashValue[163],en_end[163]);
H h164(clk,reset,0,h1InSeedSet[164],0,Hstart[164],restart[164],groupNum,hashValue[164],en_end[164]);
H h165(clk,reset,0,h1InSeedSet[165],0,Hstart[165],restart[165],groupNum,hashValue[165],en_end[165]);
H h166(clk,reset,0,h1InSeedSet[166],0,Hstart[166],restart[166],groupNum,hashValue[166],en_end[166]);
H h167(clk,reset,0,h1InSeedSet[167],0,Hstart[167],restart[167],groupNum,hashValue[167],en_end[167]);
H h168(clk,reset,0,h1InSeedSet[168],0,Hstart[168],restart[168],groupNum,hashValue[168],en_end[168]);
H h169(clk,reset,0,h1InSeedSet[169],0,Hstart[169],restart[169],groupNum,hashValue[169],en_end[169]);
H h170(clk,reset,0,h1InSeedSet[170],0,Hstart[170],restart[170],groupNum,hashValue[170],en_end[170]);
H h171(clk,reset,0,h1InSeedSet[171],0,Hstart[171],restart[171],groupNum,hashValue[171],en_end[171]);
H h172(clk,reset,0,h1InSeedSet[172],0,Hstart[172],restart[172],groupNum,hashValue[172],en_end[172]);
H h173(clk,reset,0,h1InSeedSet[173],0,Hstart[173],restart[173],groupNum,hashValue[173],en_end[173]);
H h174(clk,reset,0,h1InSeedSet[174],0,Hstart[174],restart[174],groupNum,hashValue[174],en_end[174]);
H h175(clk,reset,0,h1InSeedSet[175],0,Hstart[175],restart[175],groupNum,hashValue[175],en_end[175]);
H h176(clk,reset,0,h1InSeedSet[176],0,Hstart[176],restart[176],groupNum,hashValue[176],en_end[176]);
H h177(clk,reset,0,h1InSeedSet[177],0,Hstart[177],restart[177],groupNum,hashValue[177],en_end[177]);
H h178(clk,reset,0,h1InSeedSet[178],0,Hstart[178],restart[178],groupNum,hashValue[178],en_end[178]);
H h179(clk,reset,0,h1InSeedSet[179],0,Hstart[179],restart[179],groupNum,hashValue[179],en_end[179]);
H h180(clk,reset,0,h1InSeedSet[180],0,Hstart[180],restart[180],groupNum,hashValue[180],en_end[180]);
H h181(clk,reset,0,h1InSeedSet[181],0,Hstart[181],restart[181],groupNum,hashValue[181],en_end[181]);
H h182(clk,reset,0,h1InSeedSet[182],0,Hstart[182],restart[182],groupNum,hashValue[182],en_end[182]);
H h183(clk,reset,0,h1InSeedSet[183],0,Hstart[183],restart[183],groupNum,hashValue[183],en_end[183]);
H h184(clk,reset,0,h1InSeedSet[184],0,Hstart[184],restart[184],groupNum,hashValue[184],en_end[184]);
H h185(clk,reset,0,h1InSeedSet[185],0,Hstart[185],restart[185],groupNum,hashValue[185],en_end[185]);
H h186(clk,reset,0,h1InSeedSet[186],0,Hstart[186],restart[186],groupNum,hashValue[186],en_end[186]);
H h187(clk,reset,0,h1InSeedSet[187],0,Hstart[187],restart[187],groupNum,hashValue[187],en_end[187]);
H h188(clk,reset,0,h1InSeedSet[188],0,Hstart[188],restart[188],groupNum,hashValue[188],en_end[188]);
H h189(clk,reset,0,h1InSeedSet[189],0,Hstart[189],restart[189],groupNum,hashValue[189],en_end[189]);
H h190(clk,reset,0,h1InSeedSet[190],0,Hstart[190],restart[190],groupNum,hashValue[190],en_end[190]);
H h191(clk,reset,0,h1InSeedSet[191],0,Hstart[191],restart[191],groupNum,hashValue[191],en_end[191]);
H h192(clk,reset,0,h1InSeedSet[192],0,Hstart[192],restart[192],groupNum,hashValue[192],en_end[192]);
H h193(clk,reset,0,h1InSeedSet[193],0,Hstart[193],restart[193],groupNum,hashValue[193],en_end[193]);
H h194(clk,reset,0,h1InSeedSet[194],0,Hstart[194],restart[194],groupNum,hashValue[194],en_end[194]);
H h195(clk,reset,0,h1InSeedSet[195],0,Hstart[195],restart[195],groupNum,hashValue[195],en_end[195]);
H h196(clk,reset,0,h1InSeedSet[196],0,Hstart[196],restart[196],groupNum,hashValue[196],en_end[196]);
H h197(clk,reset,0,h1InSeedSet[197],0,Hstart[197],restart[197],groupNum,hashValue[197],en_end[197]);
H h198(clk,reset,0,h1InSeedSet[198],0,Hstart[198],restart[198],groupNum,hashValue[198],en_end[198]);
H h199(clk,reset,0,h1InSeedSet[199],0,Hstart[199],restart[199],groupNum,hashValue[199],en_end[199]);
H h200(clk,reset,0,h1InSeedSet[200],0,Hstart[200],restart[200],groupNum,hashValue[200],en_end[200]);
H h201(clk,reset,0,h1InSeedSet[201],0,Hstart[201],restart[201],groupNum,hashValue[201],en_end[201]);
H h202(clk,reset,0,h1InSeedSet[202],0,Hstart[202],restart[202],groupNum,hashValue[202],en_end[202]);
H h203(clk,reset,0,h1InSeedSet[203],0,Hstart[203],restart[203],groupNum,hashValue[203],en_end[203]);
H h204(clk,reset,0,h1InSeedSet[204],0,Hstart[204],restart[204],groupNum,hashValue[204],en_end[204]);
H h205(clk,reset,0,h1InSeedSet[205],0,Hstart[205],restart[205],groupNum,hashValue[205],en_end[205]);
H h206(clk,reset,0,h1InSeedSet[206],0,Hstart[206],restart[206],groupNum,hashValue[206],en_end[206]);
H h207(clk,reset,0,h1InSeedSet[207],0,Hstart[207],restart[207],groupNum,hashValue[207],en_end[207]);
H h208(clk,reset,0,h1InSeedSet[208],0,Hstart[208],restart[208],groupNum,hashValue[208],en_end[208]);
H h209(clk,reset,0,h1InSeedSet[209],0,Hstart[209],restart[209],groupNum,hashValue[209],en_end[209]);
H h210(clk,reset,0,h1InSeedSet[210],0,Hstart[210],restart[210],groupNum,hashValue[210],en_end[210]);
H h211(clk,reset,0,h1InSeedSet[211],0,Hstart[211],restart[211],groupNum,hashValue[211],en_end[211]);
H h212(clk,reset,0,h1InSeedSet[212],0,Hstart[212],restart[212],groupNum,hashValue[212],en_end[212]);
H h213(clk,reset,0,h1InSeedSet[213],0,Hstart[213],restart[213],groupNum,hashValue[213],en_end[213]);
H h214(clk,reset,0,h1InSeedSet[214],0,Hstart[214],restart[214],groupNum,hashValue[214],en_end[214]);
H h215(clk,reset,0,h1InSeedSet[215],0,Hstart[215],restart[215],groupNum,hashValue[215],en_end[215]);
H h216(clk,reset,0,h1InSeedSet[216],0,Hstart[216],restart[216],groupNum,hashValue[216],en_end[216]);
H h217(clk,reset,0,h1InSeedSet[217],0,Hstart[217],restart[217],groupNum,hashValue[217],en_end[217]);
H h218(clk,reset,0,h1InSeedSet[218],0,Hstart[218],restart[218],groupNum,hashValue[218],en_end[218]);
H h219(clk,reset,0,h1InSeedSet[219],0,Hstart[219],restart[219],groupNum,hashValue[219],en_end[219]);
H h220(clk,reset,0,h1InSeedSet[220],0,Hstart[220],restart[220],groupNum,hashValue[220],en_end[220]);
H h221(clk,reset,0,h1InSeedSet[221],0,Hstart[221],restart[221],groupNum,hashValue[221],en_end[221]);
H h222(clk,reset,0,h1InSeedSet[222],0,Hstart[222],restart[222],groupNum,hashValue[222],en_end[222]);
H h223(clk,reset,0,h1InSeedSet[223],0,Hstart[223],restart[223],groupNum,hashValue[223],en_end[223]);
H h224(clk,reset,0,h1InSeedSet[224],0,Hstart[224],restart[224],groupNum,hashValue[224],en_end[224]);
H h225(clk,reset,0,h1InSeedSet[225],0,Hstart[225],restart[225],groupNum,hashValue[225],en_end[225]);
H h226(clk,reset,0,h1InSeedSet[226],0,Hstart[226],restart[226],groupNum,hashValue[226],en_end[226]);
H h227(clk,reset,0,h1InSeedSet[227],0,Hstart[227],restart[227],groupNum,hashValue[227],en_end[227]);
H h228(clk,reset,0,h1InSeedSet[228],0,Hstart[228],restart[228],groupNum,hashValue[228],en_end[228]);
H h229(clk,reset,0,h1InSeedSet[229],0,Hstart[229],restart[229],groupNum,hashValue[229],en_end[229]);
H h230(clk,reset,0,h1InSeedSet[230],0,Hstart[230],restart[230],groupNum,hashValue[230],en_end[230]);
H h231(clk,reset,0,h1InSeedSet[231],0,Hstart[231],restart[231],groupNum,hashValue[231],en_end[231]);
H h232(clk,reset,0,h1InSeedSet[232],0,Hstart[232],restart[232],groupNum,hashValue[232],en_end[232]);
H h233(clk,reset,0,h1InSeedSet[233],0,Hstart[233],restart[233],groupNum,hashValue[233],en_end[233]);
H h234(clk,reset,0,h1InSeedSet[234],0,Hstart[234],restart[234],groupNum,hashValue[234],en_end[234]);
H h235(clk,reset,0,h1InSeedSet[235],0,Hstart[235],restart[235],groupNum,hashValue[235],en_end[235]);
H h236(clk,reset,0,h1InSeedSet[236],0,Hstart[236],restart[236],groupNum,hashValue[236],en_end[236]);
H h237(clk,reset,0,h1InSeedSet[237],0,Hstart[237],restart[237],groupNum,hashValue[237],en_end[237]);
H h238(clk,reset,0,h1InSeedSet[238],0,Hstart[238],restart[238],groupNum,hashValue[238],en_end[238]);
H h239(clk,reset,0,h1InSeedSet[239],0,Hstart[239],restart[239],groupNum,hashValue[239],en_end[239]);
H h240(clk,reset,0,h1InSeedSet[240],0,Hstart[240],restart[240],groupNum,hashValue[240],en_end[240]);
H h241(clk,reset,0,h1InSeedSet[241],0,Hstart[241],restart[241],groupNum,hashValue[241],en_end[241]);
H h242(clk,reset,0,h1InSeedSet[242],0,Hstart[242],restart[242],groupNum,hashValue[242],en_end[242]);
H h243(clk,reset,0,h1InSeedSet[243],0,Hstart[243],restart[243],groupNum,hashValue[243],en_end[243]);
H h244(clk,reset,0,h1InSeedSet[244],0,Hstart[244],restart[244],groupNum,hashValue[244],en_end[244]);
H h245(clk,reset,0,h1InSeedSet[245],0,Hstart[245],restart[245],groupNum,hashValue[245],en_end[245]);
H h246(clk,reset,0,h1InSeedSet[246],0,Hstart[246],restart[246],groupNum,hashValue[246],en_end[246]);
H h247(clk,reset,0,h1InSeedSet[247],0,Hstart[247],restart[247],groupNum,hashValue[247],en_end[247]);
H h248(clk,reset,0,h1InSeedSet[248],0,Hstart[248],restart[248],groupNum,hashValue[248],en_end[248]);
H h249(clk,reset,0,h1InSeedSet[249],0,Hstart[249],restart[249],groupNum,hashValue[249],en_end[249]);
H h250(clk,reset,0,h1InSeedSet[250],0,Hstart[250],restart[250],groupNum,hashValue[250],en_end[250]);
H h251(clk,reset,0,h1InSeedSet[251],0,Hstart[251],restart[251],groupNum,hashValue[251],en_end[251]);
H h252(clk,reset,0,h1InSeedSet[252],0,Hstart[252],restart[252],groupNum,hashValue[252],en_end[252]);
H h253(clk,reset,0,h1InSeedSet[253],0,Hstart[253],restart[253],groupNum,hashValue[253],en_end[253]);
H h254(clk,reset,0,h1InSeedSet[254],0,Hstart[254],restart[254],groupNum,hashValue[254],en_end[254]);
H h255(clk,reset,0,h1InSeedSet[255],0,Hstart[255],restart[255],groupNum,hashValue[255],en_end[255]);
H h256(clk,reset,0,h1InSeedSet[256],0,Hstart[256],restart[256],groupNum,hashValue[256],en_end[256]);
H h257(clk,reset,0,h1InSeedSet[257],0,Hstart[257],restart[257],groupNum,hashValue[257],en_end[257]);
H h258(clk,reset,0,h1InSeedSet[258],0,Hstart[258],restart[258],groupNum,hashValue[258],en_end[258]);
H h259(clk,reset,0,h1InSeedSet[259],0,Hstart[259],restart[259],groupNum,hashValue[259],en_end[259]);
H h260(clk,reset,0,h1InSeedSet[260],0,Hstart[260],restart[260],groupNum,hashValue[260],en_end[260]);
H h261(clk,reset,0,h1InSeedSet[261],0,Hstart[261],restart[261],groupNum,hashValue[261],en_end[261]);
H h262(clk,reset,0,h1InSeedSet[262],0,Hstart[262],restart[262],groupNum,hashValue[262],en_end[262]);
H h263(clk,reset,0,h1InSeedSet[263],0,Hstart[263],restart[263],groupNum,hashValue[263],en_end[263]);
H h264(clk,reset,0,h1InSeedSet[264],0,Hstart[264],restart[264],groupNum,hashValue[264],en_end[264]);
H h265(clk,reset,0,h1InSeedSet[265],0,Hstart[265],restart[265],groupNum,hashValue[265],en_end[265]);
H h266(clk,reset,0,h1InSeedSet[266],0,Hstart[266],restart[266],groupNum,hashValue[266],en_end[266]);
H h267(clk,reset,0,h1InSeedSet[267],0,Hstart[267],restart[267],groupNum,hashValue[267],en_end[267]);
H h268(clk,reset,0,h1InSeedSet[268],0,Hstart[268],restart[268],groupNum,hashValue[268],en_end[268]);
H h269(clk,reset,0,h1InSeedSet[269],0,Hstart[269],restart[269],groupNum,hashValue[269],en_end[269]);
H h270(clk,reset,0,h1InSeedSet[270],0,Hstart[270],restart[270],groupNum,hashValue[270],en_end[270]);
H h271(clk,reset,0,h1InSeedSet[271],0,Hstart[271],restart[271],groupNum,hashValue[271],en_end[271]);
H h272(clk,reset,0,h1InSeedSet[272],0,Hstart[272],restart[272],groupNum,hashValue[272],en_end[272]);
H h273(clk,reset,0,h1InSeedSet[273],0,Hstart[273],restart[273],groupNum,hashValue[273],en_end[273]);
H h274(clk,reset,0,h1InSeedSet[274],0,Hstart[274],restart[274],groupNum,hashValue[274],en_end[274]);
H h275(clk,reset,0,h1InSeedSet[275],0,Hstart[275],restart[275],groupNum,hashValue[275],en_end[275]);
H h276(clk,reset,0,h1InSeedSet[276],0,Hstart[276],restart[276],groupNum,hashValue[276],en_end[276]);
H h277(clk,reset,0,h1InSeedSet[277],0,Hstart[277],restart[277],groupNum,hashValue[277],en_end[277]);
H h278(clk,reset,0,h1InSeedSet[278],0,Hstart[278],restart[278],groupNum,hashValue[278],en_end[278]);
H h279(clk,reset,0,h1InSeedSet[279],0,Hstart[279],restart[279],groupNum,hashValue[279],en_end[279]);
H h280(clk,reset,0,h1InSeedSet[280],0,Hstart[280],restart[280],groupNum,hashValue[280],en_end[280]);
H h281(clk,reset,0,h1InSeedSet[281],0,Hstart[281],restart[281],groupNum,hashValue[281],en_end[281]);
H h282(clk,reset,0,h1InSeedSet[282],0,Hstart[282],restart[282],groupNum,hashValue[282],en_end[282]);
H h283(clk,reset,0,h1InSeedSet[283],0,Hstart[283],restart[283],groupNum,hashValue[283],en_end[283]);
H h284(clk,reset,0,h1InSeedSet[284],0,Hstart[284],restart[284],groupNum,hashValue[284],en_end[284]);
H h285(clk,reset,0,h1InSeedSet[285],0,Hstart[285],restart[285],groupNum,hashValue[285],en_end[285]);
H h286(clk,reset,0,h1InSeedSet[286],0,Hstart[286],restart[286],groupNum,hashValue[286],en_end[286]);
H h287(clk,reset,0,h1InSeedSet[287],0,Hstart[287],restart[287],groupNum,hashValue[287],en_end[287]);
H h288(clk,reset,0,h1InSeedSet[288],0,Hstart[288],restart[288],groupNum,hashValue[288],en_end[288]);
H h289(clk,reset,0,h1InSeedSet[289],0,Hstart[289],restart[289],groupNum,hashValue[289],en_end[289]);
H h290(clk,reset,0,h1InSeedSet[290],0,Hstart[290],restart[290],groupNum,hashValue[290],en_end[290]);
H h291(clk,reset,0,h1InSeedSet[291],0,Hstart[291],restart[291],groupNum,hashValue[291],en_end[291]);
H h292(clk,reset,0,h1InSeedSet[292],0,Hstart[292],restart[292],groupNum,hashValue[292],en_end[292]);
H h293(clk,reset,0,h1InSeedSet[293],0,Hstart[293],restart[293],groupNum,hashValue[293],en_end[293]);
H h294(clk,reset,0,h1InSeedSet[294],0,Hstart[294],restart[294],groupNum,hashValue[294],en_end[294]);
H h295(clk,reset,0,h1InSeedSet[295],0,Hstart[295],restart[295],groupNum,hashValue[295],en_end[295]);
H h296(clk,reset,0,h1InSeedSet[296],0,Hstart[296],restart[296],groupNum,hashValue[296],en_end[296]);
H h297(clk,reset,0,h1InSeedSet[297],0,Hstart[297],restart[297],groupNum,hashValue[297],en_end[297]);
H h298(clk,reset,0,h1InSeedSet[298],0,Hstart[298],restart[298],groupNum,hashValue[298],en_end[298]);
H h299(clk,reset,0,h1InSeedSet[299],0,Hstart[299],restart[299],groupNum,hashValue[299],en_end[299]);
H h300(clk,reset,0,h1InSeedSet[300],0,Hstart[300],restart[300],groupNum,hashValue[300],en_end[300]);
endmodule