`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/04/17 10:14:36
// Design Name: 
// Module Name: mpc_simulate
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`define tapesLength 16*2295
`define msgsLength (255+3*4*85)*16
`define one_msgsLength 255+3*4*85
`define state_mask_length 255*16
module compute_whitening_key(
    input [254:0] key0,
    output [254:0] key
    );
    
    wire [254:0] and_result0;
    wire [254:0] and_result1;
    wire [254:0] and_result2;
    wire [254:0] and_result3;
    wire [254:0] and_result4;
    wire [254:0] and_result5;
    wire [254:0] and_result6;
    wire [254:0] and_result7;
    wire [254:0] and_result8;
    wire [254:0] and_result9;
    wire [254:0] and_result10;
    wire [254:0] and_result11;
    wire [254:0] and_result12;
    wire [254:0] and_result13;
    wire [254:0] and_result14;
    wire [254:0] and_result15;
    wire [254:0] and_result16;
    wire [254:0] and_result17;
    wire [254:0] and_result18;
    wire [254:0] and_result19;
    wire [254:0] and_result20;
    wire [254:0] and_result21;
    wire [254:0] and_result22;
    wire [254:0] and_result23;
    wire [254:0] and_result24;
    wire [254:0] and_result25;
    wire [254:0] and_result26;
    wire [254:0] and_result27;
    wire [254:0] and_result28;
    wire [254:0] and_result29;
    wire [254:0] and_result30;
    wire [254:0] and_result31;
    wire [254:0] and_result32;
    wire [254:0] and_result33;
    wire [254:0] and_result34;
    wire [254:0] and_result35;
    wire [254:0] and_result36;
    wire [254:0] and_result37;
    wire [254:0] and_result38;
    wire [254:0] and_result39;
    wire [254:0] and_result40;
    wire [254:0] and_result41;
    wire [254:0] and_result42;
    wire [254:0] and_result43;
    wire [254:0] and_result44;
    wire [254:0] and_result45;
    wire [254:0] and_result46;
    wire [254:0] and_result47;
    wire [254:0] and_result48;
    wire [254:0] and_result49;
    wire [254:0] and_result50;
    wire [254:0] and_result51;
    wire [254:0] and_result52;
    wire [254:0] and_result53;
    wire [254:0] and_result54;
    wire [254:0] and_result55;
    wire [254:0] and_result56;
    wire [254:0] and_result57;
    wire [254:0] and_result58;
    wire [254:0] and_result59;
    wire [254:0] and_result60;
    wire [254:0] and_result61;
    wire [254:0] and_result62;
    wire [254:0] and_result63;
    wire [254:0] and_result64;
    wire [254:0] and_result65;
    wire [254:0] and_result66;
    wire [254:0] and_result67;
    wire [254:0] and_result68;
    wire [254:0] and_result69;
    wire [254:0] and_result70;
    wire [254:0] and_result71;
    wire [254:0] and_result72;
    wire [254:0] and_result73;
    wire [254:0] and_result74;
    wire [254:0] and_result75;
    wire [254:0] and_result76;
    wire [254:0] and_result77;
    wire [254:0] and_result78;
    wire [254:0] and_result79;
    wire [254:0] and_result80;
    wire [254:0] and_result81;
    wire [254:0] and_result82;
    wire [254:0] and_result83;
    wire [254:0] and_result84;
    wire [254:0] and_result85;
    wire [254:0] and_result86;
    wire [254:0] and_result87;
    wire [254:0] and_result88;
    wire [254:0] and_result89;
    wire [254:0] and_result90;
    wire [254:0] and_result91;
    wire [254:0] and_result92;
    wire [254:0] and_result93;
    wire [254:0] and_result94;
    wire [254:0] and_result95;
    wire [254:0] and_result96;
    wire [254:0] and_result97;
    wire [254:0] and_result98;
    wire [254:0] and_result99;
    wire [254:0] and_result100;
    wire [254:0] and_result101;
    wire [254:0] and_result102;
    wire [254:0] and_result103;
    wire [254:0] and_result104;
    wire [254:0] and_result105;
    wire [254:0] and_result106;
    wire [254:0] and_result107;
    wire [254:0] and_result108;
    wire [254:0] and_result109;
    wire [254:0] and_result110;
    wire [254:0] and_result111;
    wire [254:0] and_result112;
    wire [254:0] and_result113;
    wire [254:0] and_result114;
    wire [254:0] and_result115;
    wire [254:0] and_result116;
    wire [254:0] and_result117;
    wire [254:0] and_result118;
    wire [254:0] and_result119;
    wire [254:0] and_result120;
    wire [254:0] and_result121;
    wire [254:0] and_result122;
    wire [254:0] and_result123;
    wire [254:0] and_result124;
    wire [254:0] and_result125;
    wire [254:0] and_result126;
    wire [254:0] and_result127;
    wire [254:0] and_result128;
    wire [254:0] and_result129;
    wire [254:0] and_result130;
    wire [254:0] and_result131;
    wire [254:0] and_result132;
    wire [254:0] and_result133;
    wire [254:0] and_result134;
    wire [254:0] and_result135;
    wire [254:0] and_result136;
    wire [254:0] and_result137;
    wire [254:0] and_result138;
    wire [254:0] and_result139;
    wire [254:0] and_result140;
    wire [254:0] and_result141;
    wire [254:0] and_result142;
    wire [254:0] and_result143;
    wire [254:0] and_result144;
    wire [254:0] and_result145;
    wire [254:0] and_result146;
    wire [254:0] and_result147;
    wire [254:0] and_result148;
    wire [254:0] and_result149;
    wire [254:0] and_result150;
    wire [254:0] and_result151;
    wire [254:0] and_result152;
    wire [254:0] and_result153;
    wire [254:0] and_result154;
    wire [254:0] and_result155;
    wire [254:0] and_result156;
    wire [254:0] and_result157;
    wire [254:0] and_result158;
    wire [254:0] and_result159;
    wire [254:0] and_result160;
    wire [254:0] and_result161;
    wire [254:0] and_result162;
    wire [254:0] and_result163;
    wire [254:0] and_result164;
    wire [254:0] and_result165;
    wire [254:0] and_result166;
    wire [254:0] and_result167;
    wire [254:0] and_result168;
    wire [254:0] and_result169;
    wire [254:0] and_result170;
    wire [254:0] and_result171;
    wire [254:0] and_result172;
    wire [254:0] and_result173;
    wire [254:0] and_result174;
    wire [254:0] and_result175;
    wire [254:0] and_result176;
    wire [254:0] and_result177;
    wire [254:0] and_result178;
    wire [254:0] and_result179;
    wire [254:0] and_result180;
    wire [254:0] and_result181;
    wire [254:0] and_result182;
    wire [254:0] and_result183;
    wire [254:0] and_result184;
    wire [254:0] and_result185;
    wire [254:0] and_result186;
    wire [254:0] and_result187;
    wire [254:0] and_result188;
    wire [254:0] and_result189;
    wire [254:0] and_result190;
    wire [254:0] and_result191;
    wire [254:0] and_result192;
    wire [254:0] and_result193;
    wire [254:0] and_result194;
    wire [254:0] and_result195;
    wire [254:0] and_result196;
    wire [254:0] and_result197;
    wire [254:0] and_result198;
    wire [254:0] and_result199;
    wire [254:0] and_result200;
    wire [254:0] and_result201;
    wire [254:0] and_result202;
    wire [254:0] and_result203;
    wire [254:0] and_result204;
    wire [254:0] and_result205;
    wire [254:0] and_result206;
    wire [254:0] and_result207;
    wire [254:0] and_result208;
    wire [254:0] and_result209;
    wire [254:0] and_result210;
    wire [254:0] and_result211;
    wire [254:0] and_result212;
    wire [254:0] and_result213;
    wire [254:0] and_result214;
    wire [254:0] and_result215;
    wire [254:0] and_result216;
    wire [254:0] and_result217;
    wire [254:0] and_result218;
    wire [254:0] and_result219;
    wire [254:0] and_result220;
    wire [254:0] and_result221;
    wire [254:0] and_result222;
    wire [254:0] and_result223;
    wire [254:0] and_result224;
    wire [254:0] and_result225;
    wire [254:0] and_result226;
    wire [254:0] and_result227;
    wire [254:0] and_result228;
    wire [254:0] and_result229;
    wire [254:0] and_result230;
    wire [254:0] and_result231;
    wire [254:0] and_result232;
    wire [254:0] and_result233;
    wire [254:0] and_result234;
    wire [254:0] and_result235;
    wire [254:0] and_result236;
    wire [254:0] and_result237;
    wire [254:0] and_result238;
    wire [254:0] and_result239;
    wire [254:0] and_result240;
    wire [254:0] and_result241;
    wire [254:0] and_result242;
    wire [254:0] and_result243;
    wire [254:0] and_result244;
    wire [254:0] and_result245;
    wire [254:0] and_result246;
    wire [254:0] and_result247;
    wire [254:0] and_result248;
    wire [254:0] and_result249;
    wire [254:0] and_result250;
    wire [254:0] and_result251;
    wire [254:0] and_result252;
    wire [254:0] and_result253;
    wire [254:0] and_result254;
    

assign and_result0=key0^255'b011101000001110101100101000100110111000111000100100101000100111011010001111101111111001000010000110110100111110111001010010110011111110011010010100100010011110110000010111000010001111000000001111011110101010011101000100011111110111011110010100001110100100;
assign and_result1=key0^255'b110110111000010010010110001101001001111010110010010000100001000100101000111011011011001111011101010101000011011011011000111100101110111110000111111111011000100000010010000001101011000011111110001110111110011101000101110001111100101010000001101100001010100;
assign and_result2=key0^255'b100010011001100010101001111110111001100101110010000000010011110100010110101110101110110110010001101000011000100100101010000011010101001001000000101001101011010011100001000011100110100011011100100011011101000111001010001010011011100111010001101001101100001;
assign and_result3=key0^255'b000010000100011111110101001010100101101001110100111000110100110000000111000000001011001101011111000010111000011000000101101100011001001100101110001000001011010011000001110100010110001001011110100101110101010001101110000001100111101111011000010111110000110;
assign and_result4=key0^255'b001001010101011100001111100100100110011111111001011110110001100100001110111101101000010100011110010011010001100000110000100010100110010110100110101110111101010111010111001011010011110011101101010100001011010010111011011010001010000000011101000010101111001;
assign and_result5=key0^255'b011010010011111111111010101011000001000100101000000100011100011010010110100111101011100100101101011101100011001011011110001101011010001010001101111010000100100000101011100111100001011000011011000010101111101111100001000001000100000001001000000100101111000;
assign and_result6=key0^255'b101011100011110011100101000010010000010001111011001001011010010110011001011001011001110110001100001010000010011111010011111110000100001111101001011101110010101000011110100110101100111011100000101100000001101010101111110110100110011100001011111110101101110;
assign and_result7=key0^255'b100001110100101001011111111101101111101110111010101000101111101101111001111110110100011010010001100000110011111011000011011000000000000111011101011001111110101000110100101111100001101011111001011001111011101011100110000101010100111011111110110001010101101;
assign and_result8=key0^255'b010000111010110000000011110011011111010001110000001010111110100011011100011011001101101010000101010001001101001101111010011100001111011110010010001110000010010001100111101111100101000101001101110111010111010111100010101100001100111001001000010011101011100;
assign and_result9=key0^255'b010011011101100000000111001100100101010111010011001110100011000111010111000011100000100101100000011110011101001010101011000000100111110000100110110110000111001000001001100010010111111001000101000001111111111001001000000001110111101111110111010110010000001;
assign and_result10=key0^255'b100100001101110001111110001111110011011111010011111100111010010011101110100000010110100011110111101001001110011010011010001000111100110011100011101111001011111111100100111000100011101111111010001110010001110010000111010100110101011110100110100111010101100;
assign and_result11=key0^255'b100100011111000001100111011100001101011011110111011010000110000110000101010011010011010010000000001100001000001001000101011001100000011010100011011011101100000011001010010100001011011010101010100011010111011110100000100010000110010001010000010110010101000;
assign and_result12=key0^255'b000100011010010011001001000100000011010011011111010010101001011100001101110010110101001011101000010110011011000100111100110011111010111111000001100100000111110101001011000010011010111100011111000101000111001001000111111111101110011001011110011100101011101;
assign and_result13=key0^255'b101100010111100110100110100011010110000000011101111010000001001000100001000010001110111000010110111110001101111001000011101111100001110010001110110001010111000011100101010001000110000011111010011000010000100001011110101111100100011111100011000101111100110;
assign and_result14=key0^255'b100100110000001110000100110110101100011000110000100001010011011110000101011000010111001011000111011011111101100001001110000010110110111101000001011111010110010010111110000001111000000100000001000001101001100010111000100101101000001000001000000111100101000;
assign and_result15=key0^255'b101000100000100101011011010110001001001111011101111111101011010110100010000101000101100010100101001100101101110001100010001000001111100001010100001000001001101010010101000110100011001001010100001100000110111100011110110111011001010001111110111011100010101;
assign and_result16=key0^255'b110111000010000101011110011011100000011101000010000100100001100010111011011010001010111111101010001011111010101000100001001110001010110010111001011000110110111000001000110000101101010110101001011100100100110000010100011101101110001111011111000001010100011;
assign and_result17=key0^255'b001101010111101110000101110011111001111111010111111000000101001110100010110000110100111110000001111100001111100100011010000011010011100100000000101100010001100100111110110100010001010101001101011100010110101111110100001011110010011000101110100100001111011;
assign and_result18=key0^255'b100000110001000010110011101011110000111100111110000001000110100010111001110001011101100010100110010010101011110101000110110101101110111000010111000000010011100010101000000001000100101000110110111000001011011000111001111101001001110100101101010001111111110;
assign and_result19=key0^255'b110111110101100100100001100010010011101111110011000101010000101101011010011101110011000111000010010001110010010101101010000010111011010110100011011100110110101111011100000100001000011010001111100010110110100111011010101000100100110010011001110000001100110;
assign and_result20=key0^255'b101011011000101011100010110010011000010100101111110110100001000011001101001111111101010101111010000110111100101000101001101001001010111110011111011101001110100110101101100011100001101101100001101011010001010100110000000110010001101010100100101000101010110;
assign and_result21=key0^255'b000111000111111101001000110011000111100001001001011111101011100011011011111110110001011011100100000000001100110100010101111110101110111100010110101110110101111101110001000101100011100101101111010111001011100110011010101110010111011011101101010001111001000;
assign and_result22=key0^255'b000111110000110101001011000111011111111001110011111001011110011111000111001101100011001010100011001100100010101101011001110111011100101110010011100010100111100110101110001010011100000110000010010010111010100000110001111111111000111111111100001000010100000;
assign and_result23=key0^255'b001101100101101000001101010111011000000010101010111110001011111100101010101100000111101110100111110010111011011101100101000001001101111100111111000000001101000111011100010110111110010000000100110011110011011000001010110001010100011011101001110000110111000;
assign and_result24=key0^255'b010101010110100100111010100101000101101011111101101111010100111011010011011010001101111101011010001010011001011111000001110011010100001000100001110111111110010000001011100000001001001001101001111000011100011001110010011101110110110111001110100001101010000;
assign and_result25=key0^255'b000101110011011011011100101001111101011011011010101001101001010101000010100011010101000011000000111000010101011101011111110010010011111001100010110100101100011010110001100010110110010011010010010010101010100001000110001001100111101111001100101111101000001;
assign and_result26=key0^255'b101001001001100001011010010100011000001110100000111101000001100010110010110110001111001000111100100100001111111001110101110101011001001000001000101001110001100010010001101111111000000111101011111010011111000010100001011010011101000100100000010100100010101;
assign and_result27=key0^255'b010011100011011000110001000110000000001111100110100100001101101010000001000100010011010011001110011011100111111100010110001000001111011110111111011011010011010101000010101010100010111011011011001111011011101000101101110110000100001100111111100101111111110;
assign and_result28=key0^255'b011001110101010111001111010100101111101011100011010111100111011010000011101100111011001011010111110010011011111010010000000000010000100010000101001110101101000000011011001111010110010010000001100001001111100111101000010100100000001000011110111001111110000;
assign and_result29=key0^255'b110001000000011000110001011000011000001011100001111001010010000100001010000001001111110001100011011001001110111111001111000100000100100111001101001111111111010100011101101110010111110000110101110001100110101100000001111000001101110111100011100111000100101;
assign and_result30=key0^255'b011001000101011000110001111100100011101110100011000101110101010001001100111011000101111111110110100111010110010001111010110111101011011111010110010010110110010100101001000010111101001000111100011011001000000011000100110100100011111010100010111110101000111;
assign and_result31=key0^255'b110010000000000010010001011110110110010110011000001010111000100000110011100001111110000100110000000010110100001111100101000110110001010000011111010101100001110100000000101111000001111000011001101010100011101011001001000001100111001010110111101000101010000;   
assign and_result32=key0^255'b000011111011110001010010100011100110000000000110000011010000101111010101010100001111101100101011000101001010111101111110001100101001001110000011101100010100010101011000110111010011001000111011001110100011100010111101101010110010000001000001010011011101011;   
assign and_result33=key0^255'b010110100100111111100110111001111101101000100000111011000001110111100110000100010000100110010010000110001000101100111111010100110011100010111110111011010101000011000010010001101011001000000100101010000100000100111010101111111111011001001111110100111110100;   
assign and_result34=key0^255'b011011000111101001011011011111110000101010100011001100000101011101001000100110011101010110000110011001010101000111010110101000111001011111001001110110010000010011000111000111000001111110101100001100000101000110011011110011010001001101000010010010111101100;   
assign and_result35=key0^255'b111101110000111000101000000100100001111110101101010001110101111011100011110001010001100111000000101110111100101010001101111001110010111111001100100110111010001110100111110101000101000111100100010010100101010000000001010011010011000010110111111000110101011;   
assign and_result36=key0^255'b100010111111001101101010101110011101100100111001000011010111111111001010101100101111110110011001110000010111101110111011111101100000011001001100111000100000110011100000011100010010100110100010001010101100001000000011001011110011011100010110000011100001011;   
assign and_result37=key0^255'b111100000110111100010101111111101000111010010001000001111010001011110101010111100001110011100100101101000110001111101110011001111101111111000010111001111001001100110101011010101110111001010000100111101011010011101000101100011111100011100000011110100010111;   
assign and_result38=key0^255'b011100010111100110111110001001100110111101000111110100001101011100110111010100011001110010110010101100000101110100011111010011010101100111100001111101011000000111110011101101001011011011010101101010111000101010101101111010000100100100111111010010000110111;   
assign and_result39=key0^255'b001010001101001111111010000000001010010001101011010010011000111000011011111111100100011100110011111000010011111011101110000111110001101011101011101010110110110101001100000111011101101101010010010100010111101110111000011001000011110100000100011010111000010;   
assign and_result40=key0^255'b110110010101100101000100110000110101110101111110111111111000010000010011101100101101000001001010010101111101101000000101000010010101100101000011100000001011010111111010010100000001011100001011001101100101100101100001101011100011101011001010111111001110010;   
assign and_result41=key0^255'b001001000100010000110110001000100110010011011010101100100110010010101111101010100111101110000110000001010001100110010001101001011111101000011110000110100000110101101110010000101101011011100010000010010111110110010000001000000001010111011000001011101000111;   
assign and_result42=key0^255'b110011100111001111100111000000111000000011000111001000101100010110101000111100000101010000101000001001111110010111110110001010010110011101011110011001001111101000010010100001101000100110111100101001110110011010110111000001111010000100010110100011001111101;   
assign and_result43=key0^255'b100100011111010100101110101010010011001010010101110010101011011000111011000001100011001010100101000000101001000010111100011110101000111000000100000100000000011110101110000110000010010001011010011100001001011100100001111111100001100001111110000101011010110;   
assign and_result44=key0^255'b000101110000100011110111111001011011001110110111100110101011000001110111111011101001001000100100000110110100111000100010110100111110110101100000010011001110011000110101110110001001100100011000011001111001010011011100010011110001110011110100111101110001111;   
assign and_result45=key0^255'b000101000000000000000011011100010000100011011011110111100010001000100110011110100001100011010100010001010000111101111111010001001101101001100011100111111010110010011010001100011010110011110100111110001110000010111000110111010001111100010100100110111111110;   
assign and_result46=key0^255'b000101100011110010101000010111111000001101001011001110101111010010101110100111010111110011001100111011010001000011100001100010011100111101010011110001000101001111001110100011110110100000111101010001011001101111010110010101101010101011001100010001110001000;   
assign and_result47=key0^255'b000011101000111011011111110011000010110000001001100100101011001001111001111100111011011000101110001111110110111100110010010101010101001010101111011111111110010100011111011101001011001100100001110101110011100110010010101000010100000011001001111100111001100;   
assign and_result48=key0^255'b011111110111000110000101011111101011100110101110000011010101011001111101010100101101101100010100111011101000011110110001010011010000010001010100111011101111101000010010000010010110000011010110110000100011000100111100011011101001110001000000011111100001010;   
assign and_result49=key0^255'b011100011101101100110110101110110111010010111000011011000001101100011110111110011101111110000011111100001000111101010101111101000011011100000110100010101111101100100011110100000110011000000100111001111101001000110001110100100101010101110011100010011001010;   
assign and_result50=key0^255'b001100110001100001100101100111000101001111010010010010001111000010001100010001111010011001010111000101101011010101111111110000001110010001111001101100100001000110000110110011111001010001100110000010001101001011000110100111110111000010100001001001101110100;   
assign and_result51=key0^255'b011111011010111010101101001110011000111101101011111101010110100100000010100110111110101110100100100001111111101000111001001101010000101001010111001111111100010011011001011111010001010001111001111000011100111111101000100001011010011010111000110100101000001;   
assign and_result52=key0^255'b001101101100010101000010011111000110001100110010010100000111011010111001010010100011000101011011000101010001101011001101111101010010010100100001100000010111100110011011001101110111101001110101010001111100011100101101111001110100100110010100101101101101101;   
assign and_result53=key0^255'b011010101101110101111010100100010011101000011101101100111100100101011000010011111000011111110100001001101010110000101111110111110100101010101101011111001011100100111101011011100111001101110101001100110110000100111111000100011101111110001011111101011100011;   
assign and_result54=key0^255'b111010100101111100100011001010101000010011111100000010101001110100111110100000101101101101101100001001000011111111011101011000001011011011000101110010111110100011010011011011110101000101011100000111011100010001001100000110011100001101101000010111101010011;   
assign and_result55=key0^255'b111011001110111110010111101101000011001110101100001001001010011110001010101000011110100101000010000010011111110100111000000011010001101100110000110011110110100011111101000100001101100001101101011001000000011011010001101010100010011010101000101011110011101;   
assign and_result56=key0^255'b001110101101100010111111011100101000010011011001010011111101110101010100100001000101000100010111000100100010100001110110001001110100101011000111010010011110001111001001000100110101111110110100000101001110111110100001010100110101101010001010100100000011100;   
assign and_result57=key0^255'b010101110100010110001100010100111011110001101101111110101011010001011101100111111000001111100010000100101110111011000110001010101101111011111100011100000001010011011100101100010000001111010001001111001100100110000110110100001101000100010011011111111101011;   
assign and_result58=key0^255'b010100011101000010110001101111111011111111100001100000100001001011011011110010111111011110011101100110100100111111001100101010110110100010001100000101000011001011010011111011011011011010001011011110011101011000001010011011111111010100000101001010010111000;   
assign and_result59=key0^255'b111010110110010011011010110001001000101101001111100011001001110011000100101111010011100100000010111011001101010100000110101011001001100111111001101101101110111011110100100000001100011101010100010001010100111100101101001110110100000001101100110111100101111;   
assign and_result60=key0^255'b010010111011001100001010111010101110011100101011110110110111110110101010111011001111110110110011011100111010111110011000100011001110001011000110111110001110010010000110111110001110001100110110010101000011101011110000001110110111011101111001011111110110010;   
assign and_result61=key0^255'b111101011011000000011110100100011011101011011001111011000100010000001111010111010011110010010100001110010011011011011101101100011111001001100010100111111001001111010110001111111101011011001101101010101011101101011110011000101010101110110010000101011000011;   
assign and_result62=key0^255'b111001000010111000101110101010110010010111000101110100111101011101000011110000111100101001001000100100110011111101111110010111000001111000110010101001010001100110000100110110000100100001000000111000111011000101110010010001111110101101101010011110111101011;   
assign and_result63=key0^255'b111000111101110110111011011001101101001001110010100000011001000001010001101010111100101001101110100011100011100011110101101000000011111110100110110011011101111011011101011110010001101110010000000000000011101011100110111110101110000101010000011100100100110;   
assign and_result64=key0^255'b100010001101011101100000001010011100011010110001110010001000100101010101110001001111000010011100101011110000100101111110000100011101110011000000010011010101010101111010110001111010010101100111010000010101000010111000110111010110101000010001100011110000101;   
assign and_result65=key0^255'b000101011110111110101001111000000110111100100011100000010110011000110111110101011010111000111100101101111111111010010101100001100010011001110011101110011101001011000001010110100110010011101100010000011000010000101011111111111100010010001110101100100100111;   
assign and_result66=key0^255'b001101010100011001100100010100110110111101101011001010101110010101011111111001010101100111001100100001101010011010110111100110110011000101000011100110101110011110010011000110010101011100101111010101100011101111000011111100100010000010101010100011010111011;   
assign and_result67=key0^255'b100100011110110101010000000010011110111011000011001011001111110010101000010010011101110010111011110101101110010110110101111100000000101001101000001000011000111011011011111101000100001110100100110000000011010101110111111010110001101101010011011010111111111;   
assign and_result68=key0^255'b110010011011101101100100010111110001100000000100110100001011100011000010111100111011111110010110001101001110101010101100000111010100101110000011011100001010000101011000110000100100101010011010101011110101001101000100000101000010011001010011100110101100111;   
assign and_result69=key0^255'b100100000011001111001111110101000111010011111010110101101100100110111011000101010110101101111001110001110110000001010001000001101010110101001100101101100110110101010000100111000101101010111001001110111010110001101110100000010011101001110011110000000010000;   
assign and_result70=key0^255'b100000011110101000000111011111010011100001101011101100100111110110101001100011110110010110110110101100101110011011110000011110110101011011001001100100100000000000011110001000111110011111001011001111011100111010000101000111111111111110111111010101111010101;   
assign and_result71=key0^255'b000110011110100000100000000001001010101110000000011001100101111010000011110111001100000011000111100100111100001000101111110010010111110011000011001011101010101010011001001001110010000001111111000000111011101100010100100110110001011101010001011111110000011;   
assign and_result72=key0^255'b111111001010000011101101001110011001001000000000110101101000111100110111101011000011011011011110000111000111110111001100010000100001001011001000001100000101001111101011011000000000000100011101001011111000111111111000111101110011001001101110101100010001111;   
assign and_result73=key0^255'b010111101110101000111001000111101001000111111010111010111110111001101010010110001000111001110100100011101010011010100000110011111011100111110011110011110101011101001101110111000110101111110010001000101100010001110010000101011100100000011111110101011011110;   
assign and_result74=key0^255'b010111010001000110101001100000111101011001011011000001100110011000001100000100000011100000001001101100000111100111010100100010011000110110110010011000111110001011011111010010000001011011010011011000010101111110010110001011000100110101011010110010101011110;   
assign and_result75=key0^255'b110101111111110000110011011010011110011010110110101101010010000000100001111011100100111000011110010110010111001110000010001010001000110010000101001101100011111011110101101111100011111000000111001100100111000111101100101011011011110001111001010101101010101;   
assign and_result76=key0^255'b111100110010100100101111001111001011101010110111111101111111000110101111111101011000010001010010100100111110111110000001111010011110001100111010100110000001101001001110010100000111100100010100010010100101010010001001001101110101100100100011110111011111010;   
assign and_result77=key0^255'b001110000111011110011111010111010111011111100111011011111110110001110111101010110110010001010101111101101111000111110010011000101100011001000100001011111000010101000100010001000100000110100011111011011110110111000000111010100111000101101101000000000110001;   
assign and_result78=key0^255'b110001110001000011111001111011011100100100100000100000100101111010101111001111100110001011001101110000111001111100110000000111000100100010000011111000010000111010011001100011111000000000000010110101010110001100101111010111010001100001010010010100111001110;   
assign and_result79=key0^255'b001110111011010011100011100101100011101111110011110010101001111011010100001010100111011101011101101001100001101101011111110001000001110111110101111000111110010011110101101011000101010011000001000011101011001111111100001101110001110111101011100011001000110;   
assign and_result80=key0^255'b000000100101011000011111001111101101100111001010100100101101110001101110111111100110110111000001101001110000111010110110111100000110101101111110010001010111001010111001100100110011100010001011111000010011101010000101111001011010000010110001011101100110000;   
assign and_result81=key0^255'b000011101110011111010011010010111000010100001111010000001111000101001111101011100111010110011001000001010100110101010100000001101011110100100001101110011011101010010100101011000110001011001010000000111110010100000110111100001111101011001100011000100000100;   
assign and_result82=key0^255'b011010011011100100010011011111111000011100000001010000110000000001000100011101110111000001001001100110010011000110010010001100110010101010111101001110110101011111111110000010000000100011010011000111001001010111000110110100111111111110011011100000100110010;   
assign and_result83=key0^255'b110001000111001111001110000001001000001000101101011001110101101101111000111011000010010000101011001011101111011100110111100110010111111111001001000001110110100000111001111101100010001000110010110110010110101010011101000000100000000010110000010010111101000;   
assign and_result84=key0^255'b101011010010100000111110111001110110111000000100111010100111100001101010100100011100110101000011100000100110001010001111001000000010110010101110011110000010101000110000101110111111001111101111100111100011110111011001011000101101011001111010010010010110010;   
assign and_result85=key0^255'b101011001101010010101001100010100001101011011101101011100000100001000000000011000011001100011100100101000001101100101100111110110011000000110010011100010110010110100100001010100011010100110111101011001101110111001011011101110110111000001100100111001111010;   
assign and_result86=key0^255'b101010111000010101101001000001010000110010011001110101101010110111011000000111100100010110000110010100010001011111101000111000000100110001010010111100111111001001010100000111001101000010010111010111001001010101000000101010110111010100100010100111100111001;   
assign and_result87=key0^255'b010111000000110011000000111100110001001011110011111011001101111100011100110100100011011010001100000100111000100001000111110000100100100111010110010011001101010011001011111010110001000010011011101110000111000100110111011001110100100111000010011100110100000;   
assign and_result88=key0^255'b001001110110101010000011000101111111101100111011011011101010101100010011001101001110010111011010011010010011100010100101100010010101010011001101011110100100110000100001110001000110010011110000010100011001010100101111100001110001010000001100101001001100010;   
assign and_result89=key0^255'b011011001111100111001111011100011111001001101000000000100000001110001111010100101011001001110101000011110110010100111100010010011101011011100010101100111110101010111100001101100011110101100110001111100011010100111110011000000101110000101001010001101000110;   
assign and_result90=key0^255'b111001111011111000100011011001101110101101001101110101011100000111001010100110011100000001011010100001001111101010011000001011110110110000011000010101000100001101000101111011111011001110000011101100110000010001011010100110101100000101101000011101110011000;   
assign and_result91=key0^255'b110101101011011101100011110011111001101010001101111000001110000001010111010001110010011101001000000101111000011001110110010111010000010111001001111101010001011010101101010001101001011101101000111100101001001101110001111000111010001101111011111101101000111;   
assign and_result92=key0^255'b000111001100100111010101111110000101011111100100100011111010100100010000111010100001111101011010000011100011110011101001010111110101011000011001111001010001010111101100110100111110001001000100000001101110100010111100101100100010111000010111011011100111110;   
assign and_result93=key0^255'b011100110100011110110011001111000010011110111001000101010011110100011010111101001011000010101110010100100011101101110000101101101100000101001010100000110111111101110110110110000011110011100100111001000011101000101011010101001111111000011100110010011100101;   
assign and_result94=key0^255'b001101010010001111111001100000110110000001110010001010010011001000111101001110101111111001110111100101111000000001011000110000101001011101001000110100110010000000110101110000100000010011101101010111110101110010110011011001111101100111001110001000100011001;   
assign and_result95=key0^255'b100010100101101100000011110100101111000101000001000101001111010010010110110110000011000111110000111110010111000010101111011111011010101010000101010000101011011101100110111100000001110001010101110100101001100000011100101011100111100001110110101101111100101;   
assign and_result96=key0^255'b101000110001111000100000010011100011110001001101101100011001110000111001000111110011100111101100001101100000110110010100001111000111111000111001000010100011100110001000001111110001110111001100100010111111011111110101000111100100011110110110111100101110000;   
assign and_result97=key0^255'b010101101111110011000100111011101110001100011000011001000010110100110011101010100111111010001110000000111010000001010011000000100000100010001000101001101111001100101101000100111111111101010111010011101000010001111110111001111100100001100010011001111111111;   
assign and_result98=key0^255'b101110100010001001101001001101101000111011100010001001011101010111110011011101100011101011101001000010110001000010100111110010000011001000000011010110010101110100111100001010001101100101011011101011110001000010101110010011111111111000101011110000001110001;   
assign and_result99=key0^255'b110111111101110100011110101011101101000010100111000011010000011100001101011011001011110000101001111000100001100110011101110011010101001001001010101011100101110010011111010000101111010001110111110011001100110111011101001101000110101100011101000001010111000;   
assign and_result100=key0^255'b111001111000111101100110110110010001100000011001111111011101110000010100000000011011010111101010111110011111100110100010000110011100110010100111001100100100001100101101100000110011011001011000100001101111010111110100100001010010011110011100111110010100110;  
assign and_result101=key0^255'b111010011000110101111100011111010001100111110000101011101010011101001011011010001010100100110110111111000101110001011101010101010000111100110111001100101010101001100010001000011100110101011001010001101100001010101010100010100100011000111010110101011100010;  
assign and_result102=key0^255'b110110111001010110100101001001011011011111101011010100110100001100001100100001110111100010110000001011101000001100110110100101100101100000100111011011010011101010010000101001110111010111100110111010110000010001011011100011001111110101011001001000000110001;  
assign and_result103=key0^255'b100101011111001000010010111010000111110000001110011111101010101110100110100001111101110110001001101001011010010100011011100011100001010100111011110010011110110010110010111010100000101000101001010001000000100010110111000011111010010101110001000011111010001;  
assign and_result104=key0^255'b100101111110001110111111100101111111111100010110010100010110001110000001101110000010001111011110011100011100000001110111001010000110111010001110111111111000011000000111011010001101100100101110011011110101101101011001100010101000010101111001000110000000110;  
assign and_result105=key0^255'b110011110101101101001011001001110101001100010010111010011101010110100010011001110010101010011111010100100010110011111011110101000001111010100110000001000101001100010001111110110011111001111100011111000100000111100111001101011001111110001101101111011011001;  
assign and_result106=key0^255'b101111011011100011010100111110101000000011111010011001011111101101111101110100101010100101101110010100110001111100111101001100000111010101001100000011110010100110011100011011111011110101100100000101111110000100011101100011111001110100010011001101111111001;  
assign and_result107=key0^255'b010001100000100011010011100010111100101101011110110001000010010000110100001110000001001100100110101100000101111100100001100000111011100110100100011101100111100100111100001111010011010001101111011100101110100000100011000100100111111111000110111100001100010;  
assign and_result108=key0^255'b011000011100001101101100010011101101110001111110100110110110011011100101101010111111100000111011011111111111000100110010000101011001001111010010110001010000111011000110100100101000100010011111011100011000100110111001001001000001100001111100001010110110110;  
assign and_result109=key0^255'b110000110110101101100010000010011111001000001110010101011000110110101101111011100011110100010111001001001100100010011010100111111101110101101110011111110001100101011001010101110100100000011101000110010001110101110101100000011111001101000110011011100011011;  
assign and_result110=key0^255'b101111101011001000110110001000000000010111010111110001000111100110110101110001100100110000111010001100110001010110000100111110001000000000010110001010100010100110101101100111100011000010000100001111111101000010100011010110001110101000111101010001010101010;  
assign and_result111=key0^255'b001110100100010010000000111011111010101010010001101001111101010101010001110011000011110101010000011101010111010011000110000101010000100001100011111110001011101011110001101001111000111011011100110010011101011100011111010011001001100001111011001100100011101;  
assign and_result112=key0^255'b001111101010110000101111101001111000001010011101001010001011111000011010110001000010000100001100100000001011010100010010010001001110100001010111011001000100011010101110101001001110010110010101101100101101010000011001011010011111111101111110010110000111101;  
assign and_result113=key0^255'b010110001001110101001000000111010100010010101110000000100000110110100100011010000010110110000111110111011111000010101011001011011001010110000111000001001000011000110101110111111010010110010100011011110010111011001100101101101000001110011111110110111010101;  
assign and_result114=key0^255'b001001110110111011011100110011000110010010111001011111111110001000111101001101011110001000000100101011010010011001011010000011100111110001100010010011010111100000001100000100001011101011100000000110111011100110011001110100000111010001000011000011101001110;  
assign and_result115=key0^255'b010101100100111001011000111001100101111010001100000000010000001110010101010011111101100010000110100100101100001100010000001000101011100101111110101011000110001111100101001111110000101010011011010110001010111100000100011000101011001000101000110001101001000;  
assign and_result116=key0^255'b000111001100101111111001011111100000011111011010100000100101000101110100111010011011011101000100011111010111010100010011001011101101000000100000110111111010001101010000010000110100101001100111000100101001000111100001111110100011100011011110100110010011111;  
assign and_result117=key0^255'b010011111100001010011001010010101101110100111100101111110000011000101001010100001011000100001000001110110101100001100100011111000010010110111011011011010011100001011111001111101101110111101110101010000011010011100111001100100010010111100110001100010001000;  
assign and_result118=key0^255'b011010001110011100010000000100100011010001000000011110001001000110011001011001001010111110011110010011101100000100100011010011110101101001101111010110000100010101100111011111101111000000001110100000110110011001111100011011110110100101001011000101110100100;  
assign and_result119=key0^255'b111111010101111101010101000010101011111110111001101000010010111110100001000101110110001101010001100101010010010011111110001000111111110000101100000001010101011001000001101010011101100000010110101101011000001001101110101010100100011000100100100010001000010;  
assign and_result120=key0^255'b011000000010111010111010101010100111011100001001000000011001110010000010110010100000001111000001101001111101010110011100010010101001101100001100101000111101000101111111000100001110001111001111100011011111000101111011100101101010110101111110101011000100111;  
assign and_result121=key0^255'b001111010010101101001010111000111101011110001010011111001111000011101011111101010000000110111100101110011100010011000001001100101000111000101011011111000101111011000100010001000000010001000100001111001011110101110101110101101011000010000111011001100100110;  
assign and_result122=key0^255'b011110100111101011111000000000001010101111111110100110011001001010100001001010111001010111001001100110101110101110111011001111101101010101101000011111100101110111001110010001111101001010001110101111011111000100100001101010000011100001110010000010001111100;  
assign and_result123=key0^255'b110111000000001011000001110001010101101101011110010101110101100100111111110100111000000110110101001001100111100000111101100100111111001110110110000110001010010111010000110110000010001001111001000110011000001011111100100001101000000011001010101011011011110;  
assign and_result124=key0^255'b000110110001011100001010100010111110000001010010100110100101001011000010110000101011110110000110001010110110001000011010110001011010110011011011100101101011101111000010110011100110011000010111110011001100111110001101000101100000100011100011101001110001010;  
assign and_result125=key0^255'b001100010001011000000100001101101101101010010011110011101001010111011000010101010110000000101101101000100110100100001100011010100101110111010110111101010001001111010000100000110011011010111000010010000101011111100111110100010110111010100101111111101011000;  
assign and_result126=key0^255'b100000011111110000111011111101001000011011011110101000001010010101010000101000111101000100010101110111101010110101010010011101110101101000000110010100110001001100001000010001010000010111100101111000010010000000000111110110011100001001000101111001110111110;  
assign and_result127=key0^255'b100010100010000011110000010100111101000011000110001101011100111011110011011101010100011010001100110111001010010111110011000000100001100101100101010101001110100111101111000010111101100100101111110110010110000110010011100001000110101111110010000010100001111;  
assign and_result128=key0^255'b010100111100000011111011001100010111100100011001111010100001011110000001100000001000001001010101010011010110011101101100111010101000110110000011011000010001101110010010111110011000011001100001101001100100101000000011010000000011101011110110101100101010010;  
assign and_result129=key0^255'b101010111110100101000001011110111001011100001101100000110101111001010111111001000011011011001011100100000001101000110110010110010011111101000101011110100011101000110001000110001101000000000110111010010000001000001111001111010011011000100101110100010010101;  
assign and_result130=key0^255'b111000110001110001000011110011100001010010011100011010000000001011010011011101001011110101010110001110011111101111111100101111001000001010011001011101111110100100011110111000010001111001101001010110000100100000010011000000000010010011100001100010010110101;  
assign and_result131=key0^255'b011011001100011001110010000100111001001100010001101011010001110010000111000111110110110111111101000101101011001111110100000001111000010110110010010000010101100110100001110000001101001010011101100100101000100000010001100010010111001011110001010100000001100;  
assign and_result132=key0^255'b111010100001000101001010001110101101111110110100101001001011010110010101011001110001100001000110100110111110100011010110111110011010100111111011110010101100001110110000010110100100100011100001010100101101100001101101001011101111101000111111110000101010101;  
assign and_result133=key0^255'b011010111100000010110001001000011000110101001101111101001001101100001110101101000011111101110111010100011100111100100010111001110000010111000001101010110100011100001000000110001010100011110000110000001101011000001010110110111101101001000001000000010101001;  
assign and_result134=key0^255'b011100001111101101000111000000100011011111011100011110001110100010011111101001100011101101001101000110110101100110110110101001010101101111000000111000000001100111101101001111001100001011000001010010111101011101110001001001001100011101000010100101011110000;  
assign and_result135=key0^255'b000000110000101110011111010001101001010010011011010000011000011111010101111101000010111010110001110100100011010100101011010100011110101110100011101100111111100110000001101000000010011010011001010110001011011110010100110000001010000001100001010011001011000;  
assign and_result136=key0^255'b101111101000111110010011111011111111101111101010100110111111000001011001011110011010001001111011111001111110011111001101100010111110110011111111111111100010000001000000001000000100011111101011110000010010001101111010000001011100011110010011000000111000010;  
assign and_result137=key0^255'b111110111001101110100011010110000111110001101010110111000111100010011010100101001010010001010101101101110110101010011010110011011000000100010100110011011100010100010110111101100100000000110010001100100100110010101110101101111100101100100100000011000100010;  
assign and_result138=key0^255'b001000101111101001000110101011110000011000100001011011010001011000001001001111111011110100011010010111110010110010001100000101000010010101101100110110110010011010101111011011000010101011011101100111001011000001001000010100000110011000011101111100100110100;  
assign and_result139=key0^255'b001110011100110001000010001111110000000010110110011011011001001100000001111101011001100110000001010110010001000000001111011101010101000111110100000111111000101000100100100101011000110110011011001010000111110101000111111010001010001010010110010010101001100;  
assign and_result140=key0^255'b011010000001011111111000011000111001111100110100010011011001000000101100011101001111100110011011110010100111000111110111100101011110101010011111100001111101010011111110001000101111010000001110010111010110010100110111010010100011001001101101101101111010101;  
assign and_result141=key0^255'b001100000100001010111001010010000001010001001011100100101001010110110000001001010000011101000110110010011011110101101100110001010010111010101110011000000110010100111001000010101100111011110001010001001110001001001101100111110111101100110111101111001111011;  
assign and_result142=key0^255'b110111001010011111101111111110100111111111110000110101001000111000111111111101011000011010111001000010111110001011111011010101000000100000001101110001011110000000011100110110101000101010000000011001010001101011101011100010011111011001010110000000110101011;  
assign and_result143=key0^255'b000001011111100100101011011110010100110001101101111010110000011001001010111100001011001000010010010111000011001100000001100001111001100111000100001011000001100111000101111001001100010111011000011011001111010100100111001000101111010110100101001011011111000;  
assign and_result144=key0^255'b000011110100100100011010011110001100110010001010000111001110001100011100010011000100111000110101101101000011010011100000011011100010101000000011111011000000111100000010001101000101111111010100010010101111001010010101011011000111100101111110000100100001001;  
assign and_result145=key0^255'b111011110001111011000110111110110100000110010101111011010010000111001111010011000101011010110110100010000011011011110101001001100110111111011111100011000100100011110110010010110110011110101110011101000010000100001100000011100111111010111101101000111110111;  
assign and_result146=key0^255'b100010100101010111110100011010110101110111011101011100010101100100010000000000010001010100111110011101010001010010011000100111101010011101010000010100111111011000000111100011000111100000000111000100101001011111001110110100111111100110100100110000000010110;  
assign and_result147=key0^255'b100000101110000001101100111111011101100101010001101101101101110101001110010010001110100010011101110010100011010101111111011100000000101010100010001011100001110001011111001011100110101001110111110110111001010011100001000010011000100011011001001111011010110;  
assign and_result148=key0^255'b110100101101100001001000001001001010100010000011101000001111001110110100001111011011001110110011011110000100110000100101100011011111011111110101000001101110110000010001110100000010000110001000100101111010000010110001101001000100011110010111101010100010011;  
assign and_result149=key0^255'b001110001100010010111100110011011000000111000110000010000111011010011111100110101010111110101111001001101100001100010011011011000110100000010000011100001100110011001001100110000001110111010000111011111011010101000010111111010101111011110001111000010010100;  
assign and_result150=key0^255'b111001100011110011110111011101100101001111001100111000100010111010011001110111111010000100100010010101100111100111110010001010110110111100101110001111001000110010100111101011101111100000011101001111110110001110100000001010111001010010001011001010000111001;  
assign and_result151=key0^255'b010001011011001001000101101110011000111000100110101100010011101100101110001000011100101010110101010100011100100110111010110000000111110001101010000111011111111100011111111110010101110011010011111001100101000010110001010101110101001100000101111110101100010;  
assign and_result152=key0^255'b100111111111010001100100000110111011000110001100001000000011110101100001010000010000100101100100110101101100010111101011111011010111110001111011101111110101011011001110111011010001000011010010001000110110000101111000010101010111010001011010011100001001011;  
assign and_result153=key0^255'b010100010000011101101010001100101111110010010110111010011000010100110100000011000010010110011101011111010010111111101001111111111000010010000101100101000100111000100110111110000101100110001010011101000011101011100011010011111010101000111100101110111110011;  
assign and_result154=key0^255'b010100010110001101011010000011111100100110011110001101101000001000001101111010000000101010110101100111000001000011101100001010111100010001110111010000000000000010100101101011010100010100101011001110110011100110111000101000101011101000110110000110101100100;  
assign and_result155=key0^255'b000100000100010100000011100001110111100111110000000100000110000100111101101001011000010001100001111010000010101100011000010110110001010011100000001011011000100110011100111100110110001101101111110010011001110101011111011111101101001101011011110100111100110;  
assign and_result156=key0^255'b011110011001000110010000000000011001110100110110001100111001100000100111100000011111001101001000110000110110100011101101111011000100010100111110111011011110100010110000011011101001011000110000011000110100001011010100111100000010101101010010101111011110001;  
assign and_result157=key0^255'b100011111101001000110100101100011010111111010000010100001101100010011100001011111001011110011100001110100111101101100100010101110000011100111111000100111100001100010011000011100000100110000001100111111010101010011100011110101101100011001110110111000111100;  
assign and_result158=key0^255'b101101000110010011101001110110101010100101011110110011000111101110110111101100000001110100000111100001011110000101001001011100111001011110010011110010101001100011000101111011010100011010010001101011000100101001100101010000110010010101100011011001010100110;  
assign and_result159=key0^255'b101010001000011001111101100100100110011111110010100011001000000000110011111001000101101001001011111001010000011110110010000111110011010010000101111100011000110011111000111110011001010001101011101011011001001101111000111011010000010110110101011010100101110;  
assign and_result160=key0^255'b100011001111111010011111001101011011111011011101100010000101101110001000010000111101111000000101110111000010001001001100111100011010010111000001111011011010011000101011001101111110000100001110001001000001010100111001111111001101011110001101000110111111101;  
assign and_result161=key0^255'b111100100010100111000010101011101100111111011101100011001010011010000010110010100000010011010111100100111111101010010101100110011110010000111100000100100100111111000011100101010100000000010010010000000001001010010011010100100100101011110110100111101100101;  
assign and_result162=key0^255'b010100001000101001010010101010111011010001000011111110010110101010001101001110001001110011111001111011101100011001001010001110010000110010001000101110001001011100000101111000100010001111010001110011000010101110000001110111100000001011001100001010001001000;  
assign and_result163=key0^255'b111011010010001110010010000011000011101011111010011010001110010000100111111010010100001100110101000011111101011011100001100000111000011101100011001101111011000011110011111000101101101101001101111100011101111010111101101010111011111110100011011011101010011;  
assign and_result164=key0^255'b100010011011011001101101111100000010010000100111001001110010100110010010110100101111110010001001111100110111000111010010100001000001011101100001001110100010010100100111001010011111001010100010111011001111011110111000000001011100011011000101000111100111011;  
assign and_result165=key0^255'b010111001111111000101010000001111000010100011100000001011001010001100100010110100001111001000000010010001010010011010111000111010110000110111011110010000011011001010110011011010010000000000001111010011110011111111111000110010110010010000000111110000100111;  
assign and_result166=key0^255'b001111010101001110010000000011101111000010110100010010011000011001111101101001111101100011100011010000101010100001011111100101100001000101011100010011010000010100110111101011111111000010000001010011010111101010011101000111100100110011110110110101000000000;  
assign and_result167=key0^255'b010110111011000010011001101101110100000010101001011011110110010111000001100110110110111001100010101000110000010001010111100101100000111100001110000010100010000001101010000101111011110110001101011100100001011011001110110110000111110111011110110010111011100;  
assign and_result168=key0^255'b111101101000010100001001110111101011010101100011000011100111101101110110110011001100110001100101000100000111100100000110001001111010010010000110000001000010110011101001100001000110100100000100010110110110011111110010010101010000000000001010100011110010101;  
assign and_result169=key0^255'b000010000000010011000101111111100001011011011110001000010001111000111111001011100110111000010010110000001000000101000010011010011011111101101100010011010001001101001101010111011110100110101000001010001111101110011001011011111010100000000110001011110000110;  
assign and_result170=key0^255'b010101101001011101011110111100101101110000001101000011100110011100111011011001100111000111100101111001101010011101100110011011000110101001110011110010011110100011100111111010110100000110111011100100110010011101010011100100110100001010001111000110100100110;  
assign and_result171=key0^255'b110111110010001101001010100101000010111110110010100111010011110000110100101110111001101111100010000111101011011000011100100011011001001000110110100100101010000001100000001000100100010111000100011000001011001110001011110010111010101100010010010000000110011;  
assign and_result172=key0^255'b001000000101110110101100110001001100111001011000100100101011101011000001111100000000011100110001100111000101101110100100001000011110110110111100001100010000110000110011001111100000000000100111101110000011001000001000000111010100011011111000111111000111001;  
assign and_result173=key0^255'b100000000010100011011010010100010101001001100100101010010100110101010001110100001010000000110010111001000100000111101000111111100101100000110100011001101000001100000110000100100001101011100011110100110010111001011001110001010011100111101110000001101111011;  
assign and_result174=key0^255'b101101000111011101100111000011100011000101010000110001110111011101000010100111001000101111111010011000000111100001011010000110010000111010010010111000111010110010100011111011001101101110010000111111011110111110100011110010001000101110011110110101101010101;  
assign and_result175=key0^255'b011110111101100100000001111011100111000001010111011100011010100000010110001010000000010010110100110110101111011111110001001011011011110110110101001011001110101010110110101101111111111011110011111000010101110011001001111000011001000111100100101101101000010;  
assign and_result176=key0^255'b010111011100101010000001110101000111100100111000011101111111000110000000010001010111101101100001000000001100001001110010010001000111000101010110100101101011000010000001100000111110011100010001000101001101101100100100101011010010010111010001001101111110000;  
assign and_result177=key0^255'b010100000010011101001101010000000001001001011010000110000111110111010111011111001001010101000001010010010001111100111010010111010100100100111000001000101111110001010100010001011110101100111000110000100000010001110110001011001001011000111101010101001011110;  
assign and_result178=key0^255'b000100101000000010001100011101111001011011000100011101110100011010101110110000000101001111011111111111001100000110100110011000110010000110011010001000011011100001110010101001011100000000010111101010100001110000100000110100011000100000101100011110000000000;  
assign and_result179=key0^255'b111001110000110111001111010111111000111000100010001000110110000111101011110111011110000000001110101110110111000011000110111111110110110111001111001011000100101011111010111010001011101110001110011101001111110000101011111001111001111100000011111011100010101;  
assign and_result180=key0^255'b011100111010000111010111010100111111111110101110010001101010101100000001010011101001011100100011000110000011110010000100011011101101110101011101011110101100101011111101101001001000000001010010010111100001101111101100010001101101000110011111110111001101100;  
assign and_result181=key0^255'b110111001011010011110110011010101010111110110111100111011010000101100101001100100100001100010011110100011111111001110100001011100101000101010010000101101101000110010110101110011100001000111110000000111100101110011110011001000000110101001101110100100101001;  
assign and_result182=key0^255'b010001010110101111000011101100111100010011001110000001110101110011101010001110100010011000001011100100101100111010111010110001000010110100000001111011111001001010000111101010000000101011010110101001101110011011011011110111100011011001011110010011111111101;  
assign and_result183=key0^255'b100101011010110100001010001010100011000011010110011010011100001100100100111010101000110111001000011011010110100000010011111001110001000111011000010100000010010101101111100001100001100010011110001011100010010100011100100110011101010101111001011100001100001;  
assign and_result184=key0^255'b101110111001100110010011101001010100101100011110001110111111110101011110000101111111001011000010100100100100010011101110010000110100001111111100000111000101111010000011001110100010000010110010101010111100101101100011101000000000100011001111101000001110000;  
assign and_result185=key0^255'b001100111011000000011011000101111110011101000011100010111000100101010110010010100111101011111110100010011000111010101101110000101000111011111011010011111011010001110010111001000100101101010000010011111010100111100100000101010011010011011010101000100001110;  
assign and_result186=key0^255'b100111000010111100000001111000010001010000000000101110010100001010110101001001101110110110111101001000011110000001000010011000011111011100010000000100111111010010101110111111000100011110100001110011101101101000010001100011011011010011110110001010011110001;  
assign and_result187=key0^255'b111111100001101100010101001111000111010101111100011011111000101110101110100011001100000000111011000110011010110110101011000001111010000110110000001001111110001001101111100110111010100101001100011001101000100001000000110000000011111010010001001011001111101;  
assign and_result188=key0^255'b011111011100101100011101111111001010001010100100010000100111010110101001110000010100111000011011100111101101010101111011101011100010101001011001011000001111011100110101101000011001101011110011010001001100101100111100011000110011011000101111100011011100101;  
assign and_result189=key0^255'b011101110000001001101110110110110101001100001011000100101011001001000000101001100100110000011011011000110000001001101100001111110001000011101101100010011110100010010011010110111001011110111000011010100100110110111011000111010101001111111001001100010010100;  
assign and_result190=key0^255'b110011111000000110010001001100110110101001110100001000110011100100001100001010111001111110001001101011000111110000001010110101010000101110001101100000011111010001011110101100000101101101111100100101110010001100010111000101001100110101110000001011100100000;  
assign and_result191=key0^255'b010110001111011000101110111111111010101100010100000110011001111011011111010101100011110101100000011000101000011011111110110011110001110100000110011000100011110111100001010100111010111111010100100110010101100011101110100000011111001001000110111101011001100;  
assign and_result192=key0^255'b000101010101011011110010111010000111000110010101111010000001101111110111010101110011111001000011100000100101101011111100001011001110100101010001110011001100000100001111001110111010011011111001000110110100011100110011111000000010010001101100001000111110111;  
assign and_result193=key0^255'b010101111001110101100101010001100011110100111111010101000000000110010100100101001010001101001100110011101110011001101010001111011101010001100000111010110101111101000101000110111000000110110111011000000011111110001010010001001101100111001101101011001110101;  
assign and_result194=key0^255'b100011110011111001101101101100001011111110000011111101001101010100010011100101100100001011011101000111100101101010110000011111010110110010101100001011011011101110111001111100101001001011000101010001111110111011001101111001000111101000111100110110100111111;  
assign and_result195=key0^255'b000011001011010100101101101110011001000100011110100111100011000101011100111110110101101100101110110110001000000010100111001110010100011101100000110100111100001010011101101100000111111111110101011011000110001000101110001111111110010001110011011101001101111;  
assign and_result196=key0^255'b010010011001001111100101011010001110001111111110110101100010000011011111010101010011010111010110011111000010111111101001000101010111111010001000011101011011011101001011001000110101010100101101001010011000111001100110011011100000111010111001011110011100000;  
assign and_result197=key0^255'b110101000010110000101011001101110010111010100111100100011000001110110110110100110101000101011000101010111001100101101111000011110011110010000110011011000111100101110010100111111100010010010101100001011101010011001100110101001010011110011001010011100011010;  
assign and_result198=key0^255'b010010101000011010010110001011100111110110000111100011010010111111111101111110011111101101110110101000000010111000011100111100001111001100110000001010000111001111111110111100000001101010101001101111001100010110101000101100110101100111100011010001001011000;  
assign and_result199=key0^255'b000010001001111001010011111011010111101101010000100111010100001010001101111010001111111010110110011000101000001000110110011010101101110000000111000111101010100101101100011111011000110110011011010110001100000010110000101111000010000011000100100000111111110;  
assign and_result200=key0^255'b000001110010000111001110010111110000000001011101010010001100100001101111010110111011001100010101001000001011101001100110001110111110100101110010110010011000001111000111001000111111111000010110101110101111111011101011001001001010110101100011001110011101111;  
assign and_result201=key0^255'b011011111011011000011010101111001111010000100010011111111111100111001101110010110111000011000010011101100111000110110010101111010000000100000010110011001010011000110111111110101001101100010011110110100000011000010111100110001010011111110001001001011100001;  
assign and_result202=key0^255'b011011001000010010011000111001000000000111010110100010000110010011000001101001100000011110100101111100001110001100100101011100111110110100010100011101011100110110110001111010100111001110010111001110101101101110111110001010010011101010111101000011000101000;  
assign and_result203=key0^255'b001001010001010000001011000010111011101100011100001111011100010100000101100000010001011011010100100101111100001011011111111111101100011011011001110101011101011110000110011011100011111100101000110100011110100101000111101001100001111101010100101101101001101;  
assign and_result204=key0^255'b111100111100010101110100011011000011110000001111100001000011000111101111111010010000110010100001110000111000001010001100010011011101000001001001011111001100010011000111111000100000101100000101011001111000000111010001111100100001101000101010010001101101010;  
assign and_result205=key0^255'b101011011010101000101011101111011100101001110000101011101000110100111010010100110010110010010000011111101010101101010101101010111000110101101000100101000011000000011000010011010000101011110001100011101011101111110001000110001111111000000100110010100011000;  
assign and_result206=key0^255'b100101110000100111101101000011100100001010011111101010001100111110001001011010111100000001010011111101010011101101011001100101111000010100001001001101010111001111000101100110011101100000110110111111001111101001110101001110001101101000111101100110001100001;  
assign and_result207=key0^255'b001011000111110000111100000001100010100101101101111111010011011101001011110110010111111111011010011100010010110011101110110011011110011010000001100101111101011000110000111010111100111110110111010000100011010000100100000110010011001111111110010001110001011;  
assign and_result208=key0^255'b011010110111111010011111001100001111110111100110000010100000010111011110011110000101011010000100111010110100101100010100100100011111000100100010000011001111000110110011101000100100100111101010111100111111100110001100110010000000100100000011011001101000000;  
assign and_result209=key0^255'b101000100111110010000000110100010010100001111110100101101111010100100001100010010101000111100101001110010010001100100010011010101111101101000011001110000111100010010010111000100101101000010100110110000011111101000110101111111001100010010101101111110101110;  
assign and_result210=key0^255'b010001111010010001000010111010100011000000010110010111100001010011111001100001000110100010000011000001101001001101001100000110111000101111100001010000011111010010000110100101111010001010001000101111101101110100100111101011000100110111001000001011000101110;  
assign and_result211=key0^255'b100001111001101011011100000011011111000100101101010111111010101010000111001001011010110110101110001101100010110101100111011111001111110110110101010101010111101001101100110101110011100011000110111101101011001000000100000110001100101110011000001111101010001;  
assign and_result212=key0^255'b010110100110111110101111010010110111100101001001101011110100000000101010011011110001000011001000011010100101001111110111101101101001001110101111001111001110010100000101010100001101000011101101101011111101001011001111010011100001001100000101001000000011100;  
assign and_result213=key0^255'b111000101010011011010111001001110001011110011101010011110101001011101000111101110001000110011110100010011111000100011011011001000001111000000111101100011111110000101111000010111011000111100000000110011100101000110111011000001011101110010111000110001111000;  
assign and_result214=key0^255'b000001111010001110111010110001101010001001010110010111000101101001000110110111001001011101011111110011101000000001000011010011110001011000000011000001100001101110111111100111001101111010000011010110111111111110010011010101101110010001001010001100001111011;  
assign and_result215=key0^255'b111010101110101001100000001100101001100110011011100111110110111110101000101100100101010010100000011011000000110111001000100010010110010110100010110000011100011000001110110110110101000110011111000011001010011011110011011001110110110100000110011000010110011;  
assign and_result216=key0^255'b101111010111100100100110111001111101101000110001110100110000001000010111100101111101001011100100101000000000000011110011110001001000110001111100011010001101001000001101000100001110001101110001011111100001011011000000111111000011001000111001010011010101100;  
assign and_result217=key0^255'b101101000101011111101001010110110011100101110010000001100010000000110001100110000000111010111011101110011101110101111101110000100110100110001011001110111011001110101001100100110011010011010100000100110010111101001101000011000000010110101001100001101001111;  
assign and_result218=key0^255'b110011001101100101011010101011110010001111001101100011000000101110001000101110001101000011000100011101010000100100100110001110010001011010010100001110001110110000110001101001010101011110001000000000111001000100010111100011111100110011011100101111000010010;  
assign and_result219=key0^255'b100011000010011011000000111011101011111010101100010110001101011001111101010110111011101110011111011110010011101100111111111100010101011011010001111011111100101101110010101000000011001110110001011010010011111110111001001100110010101101000101100011000100111;  
assign and_result220=key0^255'b010011101110001000011100001101111111001010010101101011110110011111101011101111101111000111110010111000100011110101001100001100001011100111011001111000101111000111101010100001000101110010100110101011000000111111001001110111000010010101011010011010000010000;  
assign and_result221=key0^255'b101111011100100010001011011011000111010010010100110110100101101001101010010100100110111110101101011100001010010011011010000111001100001101110000010010000011100000101110100101110111110101001010101101000010000111000000111011001111110011111100011111100110000;  
assign and_result222=key0^255'b101101011101011000000100100000111101011111010100111011000111011000110010110000101110101111111111011000101111110000101000100001001100101011101101011110100001010001011011110100111001010111100110010111111011110111000001110101110000001011101100011110010101001;  
assign and_result223=key0^255'b100000111100011011000000000010101000101010000000010010111110101000110011000100100011100101011101010110101001001100010000111001000110000010101111011001010100111011110101011101011111001000001011010000100011001001110111101000011010011010101001100011101001101;  
assign and_result224=key0^255'b011101101011110010111100000111111101101000110110101001000110011100101000100000100100001111101001010110100011001101011111111010001001011100101110000111110101000000011001001101100110101000011110101110100100000100101101101101111101101110000110011101001100010;  
assign and_result225=key0^255'b010101010001000100001010100101111100111000000000001100011110001101100000011111001110011011011010110011111010100111100100011111101110010111001011001101000000000001011001100100000100100001011111011101101101110000000100111111000011110010110110110111100010010;  
assign and_result226=key0^255'b110001111000000100011010001100010101100010011110010011000111111101000110011000001101100010100101110011000010100111010110000001111111111110011111100101101001101101100001000010000100010011100001000111001011111010111110001010101100011110101100000110011111001;  
assign and_result227=key0^255'b010111011100111011011011010111101100000110111011011000111001110111100001010100000110100110010100011111001100000010111011010100101101110111000110011110101111111010011100110000000011011001101010011101111001000001010011011101101010100110010011110111011100111;  
assign and_result228=key0^255'b101111010001110011110011110001100000010110011000111101001101001110000110000010010000111011100011111100000110011010111000110101100010011101010001000010011111001100011110011101111110100000100100111110101011110001001001010111101011011001111010101111110010111;  
assign and_result229=key0^255'b111000011110000000010110100100111001101000101101111001001011001001001000010010011000100001010101011111010101010101111001101010001010110100101111110000011011001100011000001110001111011010110011111000101111010010111010111010101111011100101001100011001110010;  
assign and_result230=key0^255'b110001011100010011010000111010011000000111000111000000110010111101111000100101101110111001000101001010100110101010000001110101111101111101000000010111110100011111011000100101001011010111101000101101101001111100011111100001101111011000001110101011010100000;  
assign and_result231=key0^255'b100000101110001001101101111000111011001010000101011111000011101000100000000001011000010101011111000110110010100110101111010011111000001100011010000110101011101001001110010000011011001000110011010000000010100111010000101100100010010011011100011100100001101;  
assign and_result232=key0^255'b010111011100100010101101001001100101100000101010111110000001011001101110101011000101100101001110010010000111010110111110000000100011111001011110100101100101110100010100011100001101001100110110101110110011010001011000011110000110011110100111100111110101100;  
assign and_result233=key0^255'b111101101101101101000100000101110100011111010000100101001101011100011111101110101001111000101101011101111100010110001011111011111011101001000001101111100101011010100111001100000010111011111001100110000000011011010111010010001100100101011001001010101010111;  
assign and_result234=key0^255'b001100011010011011101111110101010010011110110010110000100010100000100001100101101010010110101010111111101110001111100110000101001110001011001100011101101111101001011110000110010111100110010111011000101101010010011100110100001110000111010100001101111011100;  
assign and_result235=key0^255'b001111111100001001011110010100100100100100111010001001000011000001110111010100010111101100001011001011011110100011011111010000100000100000100111010110111110000110000100011110101001101000111001001000111000001111011000110010011100101011111001010110111101010;  
assign and_result236=key0^255'b010101111011110000001011011101011110110001101011100010010100100011011100010101110101111110011101001011101100110101100010110010111100011101001000010010110100010001101110001111110011000001001001010110111110011111101010010000101010111111000001100100011111100;  
assign and_result237=key0^255'b001000111011000111000110110010101101011000101111001101001000110110110100110110100110100000010101010100000100101001011001011011001001011111101101100101011111101111110000111100100000000101010111001010000111000100110100010011100011001010011011101001111000000;  
assign and_result238=key0^255'b110000111101010101100000100010010011100101011000011111100111110101100100001111101101001011001000110010110111111100111010110101101101101100001011100110000101111010001101100011110100010100101001010000010110101110000001011010000100100000101011010010101100001;  
assign and_result239=key0^255'b100001001111011101001111001001110001000100101110100110011110001011101101001001000110111001110110101011001000001010100001010110101011100001101101110110101110010001110100000110000111101100110000111001010001011001100110010111111011101100001001010111110010001;  
assign and_result240=key0^255'b011000011100000101000101010110111101010011000101100100101011011101000011001100001001001000001101100101111011101001001101101001000100100110100100000101110100000100101000110001101001100010000000101101001011100100111111000100110110011100111110100010000000110;  
assign and_result241=key0^255'b101100100111011110011100000110001110100010010101001010011000001011011010110111000100111100001001110110111111011110011101001011101111011110110000000101011000110101000111010101001101011010101111011000100001110100110010110110001000000011110010110000100100111;  
assign and_result242=key0^255'b000010010111110111101000010100011100010110010101111111000001101100001000111000000010000001011000110101011010010011001100000111101000101011100000111001111101001000101101101100011011110101111000111010111010110000011000110011000000110111111110111001100010100;  
assign and_result243=key0^255'b010000111000110010011110011001111111010001100010110101011100111000010100100001001110011010111101101101011111100001001001010101001100101111010000001000001111000001001111010011100001001100101011010010001000110111010110110010011100011100111001011001111010100;  
assign and_result244=key0^255'b010011011010001100010011111010101110101110110010010011011111110111100111010001000001011011000011100011000100010101010010100100000001011011100111010000011101100110000010100111100010010100110001101111000011000111110101100101001100100100000101000000001100111;  
assign and_result245=key0^255'b000111110100000011100010111100011110100010111001101000000000111100111110011110101101000010110111000110111101100111100011111100100011111101011001000101000011000001110010111100111001001011011111010100001101010101110110110001100100010011000100111001110000110;  
assign and_result246=key0^255'b000011111011010101110100011010111110001101010010110001011011111010110001111000110001101110001101110101010101010001011100100110110100010001101001110001010111001011100111011100110011110110011011010001010010001010001100001010110111111110000010110110001010000;  
assign and_result247=key0^255'b100001001010000101100011010100100011100000010001110101010011010100000110001111110011101011111011100001001001010010010010111010010000110110000000010001001001011001111011000111110100011100000111010101100110101010101000011111110011000110001000100011111110111;  
assign and_result248=key0^255'b010001110010111100101001001001111001011000000001100001000100001110001111100100001001001011110111001000111110010101011001001001011101110011100001010101100000101110100010001111100101001101011000000110000111111101101101001111011110000001110001010111100110001;  
assign and_result249=key0^255'b010101011011010101101111100010010111100011001010101101101101001001000010111001010101111111000101000010110010110000010011001101110101000110111000110000101101110110000111011111010010011111011111000010101101000111000001110101000000010110111010101001111001001;  
assign and_result250=key0^255'b011001100101101010011111101101010010111101101100011101111101101101010000011110110110110100110111011101010110100010001000101101000110000110001100000000000110101010000001010001001011011010010010011111010000001010110010100011111001101110011000011101011100111;  
assign and_result251=key0^255'b111001000101000001001010010100001110010010111101001110001111011101101111110100101010001010101100101111011000101001010011100010100100100000111010100110011101111010010011111110001101010100001001001000110110111100011111000000110101011010011111101100100011001;  
assign and_result252=key0^255'b101101101011000100100110000110011000000111011111001100000011111101001000000100010011101100101111000101101000010100111111010001010000111010001000011000010010111101110000010100000100101000100110000011011011010100100101111011011010000000001110111000101110110;  
assign and_result253=key0^255'b010111110110010110100101000000010100000001101110000001011011101110000101101111111000111111001111001001101100110011111001111111001000001100101001001100010100011000011110101011110001101101100011010011101011000001011011001111010111100101101100100001010000100;  
assign and_result254=key0^255'b011101100010011100001111000001000000110110011011001110101010001010110000010110000001110100001100001001111100100111101100111001111100101100101000010100101001010111010011001001010010000011010000011010110100101100101100110010110110001101100000001111101110100;
    
assign key[0]=and_result0[0]^and_result0[1]^and_result0[2]^and_result0[3]^and_result0[4]^and_result0[5]^and_result0[6]^and_result0[7]^and_result0[8]^and_result0[9]^and_result0[10]^and_result0[11]^and_result0[12]^and_result0[13]^and_result0[14]^and_result0[15]^and_result0[16]^and_result0[17]^and_result0[18]^and_result0[19]^and_result0[20]^and_result0[21]^and_result0[22]^and_result0[23]^and_result0[24]^and_result0[25]^and_result0[26]^and_result0[27]^and_result0[28]^and_result0[29]^and_result0[30]^and_result0[31]^and_result0[32]^and_result0[33]^and_result0[34]^and_result0[35]^and_result0[36]^and_result0[37]^and_result0[38]^and_result0[39]^and_result0[40]^and_result0[41]^and_result0[42]^and_result0[43]^and_result0[44]^and_result0[45]^and_result0[46]^and_result0[47]^and_result0[48]^and_result0[49]^and_result0[50]^and_result0[51]^and_result0[52]^and_result0[53]^and_result0[54]^and_result0[55]^and_result0[56]^and_result0[57]^and_result0[58]^and_result0[59]^and_result0[60]^and_result0[61]^and_result0[62]^and_result0[63]^and_result0[64]^and_result0[65]^and_result0[66]^and_result0[67]^and_result0[68]^and_result0[69]^and_result0[70]^and_result0[71]^and_result0[72]^and_result0[73]^and_result0[74]^and_result0[75]^and_result0[76]^and_result0[77]^and_result0[78]^and_result0[79]^and_result0[80]^and_result0[81]^and_result0[82]^and_result0[83]^and_result0[84]^and_result0[85]^and_result0[86]^and_result0[87]^and_result0[88]^and_result0[89]^and_result0[90]^and_result0[91]^and_result0[92]^and_result0[93]^and_result0[94]^and_result0[95]^and_result0[96]^and_result0[97]^and_result0[98]^and_result0[99]^and_result0[100]^and_result0[101]^and_result0[102]^and_result0[103]^and_result0[104]^and_result0[105]^and_result0[106]^and_result0[107]^and_result0[108]^and_result0[109]^and_result0[110]^and_result0[111]^and_result0[112]^and_result0[113]^and_result0[114]^and_result0[115]^and_result0[116]^and_result0[117]^and_result0[118]^and_result0[119]^and_result0[120]^and_result0[121]^and_result0[122]^and_result0[123]^and_result0[124]^and_result0[125]^and_result0[126]^and_result0[127]^and_result0[128]^and_result0[129]^and_result0[130]^and_result0[131]^and_result0[132]^and_result0[133]^and_result0[134]^and_result0[135]^and_result0[136]^and_result0[137]^and_result0[138]^and_result0[139]^and_result0[140]^and_result0[141]^and_result0[142]^and_result0[143]^and_result0[144]^and_result0[145]^and_result0[146]^and_result0[147]^and_result0[148]^and_result0[149]^and_result0[150]^and_result0[151]^and_result0[152]^and_result0[153]^and_result0[154]^and_result0[155]^and_result0[156]^and_result0[157]^and_result0[158]^and_result0[159]^and_result0[160]^and_result0[161]^and_result0[162]^and_result0[163]^and_result0[164]^and_result0[165]^and_result0[166]^and_result0[167]^and_result0[168]^and_result0[169]^and_result0[170]^and_result0[171]^and_result0[172]^and_result0[173]^and_result0[174]^and_result0[175]^and_result0[176]^and_result0[177]^and_result0[178]^and_result0[179]^and_result0[180]^and_result0[181]^and_result0[182]^and_result0[183]^and_result0[184]^and_result0[185]^and_result0[186]^and_result0[187]^and_result0[188]^and_result0[189]^and_result0[190]^and_result0[191]^and_result0[192]^and_result0[193]^and_result0[194]^and_result0[195]^and_result0[196]^and_result0[197]^and_result0[198]^and_result0[199]^and_result0[200]^and_result0[201]^and_result0[202]^and_result0[203]^and_result0[204]^and_result0[205]^and_result0[206]^and_result0[207]^and_result0[208]^and_result0[209]^and_result0[210]^and_result0[211]^and_result0[212]^and_result0[213]^and_result0[214]^and_result0[215]^and_result0[216]^and_result0[217]^and_result0[218]^and_result0[219]^and_result0[220]^and_result0[221]^and_result0[222]^and_result0[223]^and_result0[224]^and_result0[225]^and_result0[226]^and_result0[227]^and_result0[228]^and_result0[229]^and_result0[230]^and_result0[231]^and_result0[232]^and_result0[233]^and_result0[234]^and_result0[235]^and_result0[236]^and_result0[237]^and_result0[238]^and_result0[239]^and_result0[240]^and_result0[241]^and_result0[242]^and_result0[243]^and_result0[244]^and_result0[245]^and_result0[246]^and_result0[247]^and_result0[248]^and_result0[249]^and_result0[250]^and_result0[251]^and_result0[252]^and_result0[253]^and_result0[254];
assign key[1]=and_result1[0]^and_result1[1]^and_result1[2]^and_result1[3]^and_result1[4]^and_result1[5]^and_result1[6]^and_result1[7]^and_result1[8]^and_result1[9]^and_result1[10]^and_result1[11]^and_result1[12]^and_result1[13]^and_result1[14]^and_result1[15]^and_result1[16]^and_result1[17]^and_result1[18]^and_result1[19]^and_result1[20]^and_result1[21]^and_result1[22]^and_result1[23]^and_result1[24]^and_result1[25]^and_result1[26]^and_result1[27]^and_result1[28]^and_result1[29]^and_result1[30]^and_result1[31]^and_result1[32]^and_result1[33]^and_result1[34]^and_result1[35]^and_result1[36]^and_result1[37]^and_result1[38]^and_result1[39]^and_result1[40]^and_result1[41]^and_result1[42]^and_result1[43]^and_result1[44]^and_result1[45]^and_result1[46]^and_result1[47]^and_result1[48]^and_result1[49]^and_result1[50]^and_result1[51]^and_result1[52]^and_result1[53]^and_result1[54]^and_result1[55]^and_result1[56]^and_result1[57]^and_result1[58]^and_result1[59]^and_result1[60]^and_result1[61]^and_result1[62]^and_result1[63]^and_result1[64]^and_result1[65]^and_result1[66]^and_result1[67]^and_result1[68]^and_result1[69]^and_result1[70]^and_result1[71]^and_result1[72]^and_result1[73]^and_result1[74]^and_result1[75]^and_result1[76]^and_result1[77]^and_result1[78]^and_result1[79]^and_result1[80]^and_result1[81]^and_result1[82]^and_result1[83]^and_result1[84]^and_result1[85]^and_result1[86]^and_result1[87]^and_result1[88]^and_result1[89]^and_result1[90]^and_result1[91]^and_result1[92]^and_result1[93]^and_result1[94]^and_result1[95]^and_result1[96]^and_result1[97]^and_result1[98]^and_result1[99]^and_result1[100]^and_result1[101]^and_result1[102]^and_result1[103]^and_result1[104]^and_result1[105]^and_result1[106]^and_result1[107]^and_result1[108]^and_result1[109]^and_result1[110]^and_result1[111]^and_result1[112]^and_result1[113]^and_result1[114]^and_result1[115]^and_result1[116]^and_result1[117]^and_result1[118]^and_result1[119]^and_result1[120]^and_result1[121]^and_result1[122]^and_result1[123]^and_result1[124]^and_result1[125]^and_result1[126]^and_result1[127]^and_result1[128]^and_result1[129]^and_result1[130]^and_result1[131]^and_result1[132]^and_result1[133]^and_result1[134]^and_result1[135]^and_result1[136]^and_result1[137]^and_result1[138]^and_result1[139]^and_result1[140]^and_result1[141]^and_result1[142]^and_result1[143]^and_result1[144]^and_result1[145]^and_result1[146]^and_result1[147]^and_result1[148]^and_result1[149]^and_result1[150]^and_result1[151]^and_result1[152]^and_result1[153]^and_result1[154]^and_result1[155]^and_result1[156]^and_result1[157]^and_result1[158]^and_result1[159]^and_result1[160]^and_result1[161]^and_result1[162]^and_result1[163]^and_result1[164]^and_result1[165]^and_result1[166]^and_result1[167]^and_result1[168]^and_result1[169]^and_result1[170]^and_result1[171]^and_result1[172]^and_result1[173]^and_result1[174]^and_result1[175]^and_result1[176]^and_result1[177]^and_result1[178]^and_result1[179]^and_result1[180]^and_result1[181]^and_result1[182]^and_result1[183]^and_result1[184]^and_result1[185]^and_result1[186]^and_result1[187]^and_result1[188]^and_result1[189]^and_result1[190]^and_result1[191]^and_result1[192]^and_result1[193]^and_result1[194]^and_result1[195]^and_result1[196]^and_result1[197]^and_result1[198]^and_result1[199]^and_result1[200]^and_result1[201]^and_result1[202]^and_result1[203]^and_result1[204]^and_result1[205]^and_result1[206]^and_result1[207]^and_result1[208]^and_result1[209]^and_result1[210]^and_result1[211]^and_result1[212]^and_result1[213]^and_result1[214]^and_result1[215]^and_result1[216]^and_result1[217]^and_result1[218]^and_result1[219]^and_result1[220]^and_result1[221]^and_result1[222]^and_result1[223]^and_result1[224]^and_result1[225]^and_result1[226]^and_result1[227]^and_result1[228]^and_result1[229]^and_result1[230]^and_result1[231]^and_result1[232]^and_result1[233]^and_result1[234]^and_result1[235]^and_result1[236]^and_result1[237]^and_result1[238]^and_result1[239]^and_result1[240]^and_result1[241]^and_result1[242]^and_result1[243]^and_result1[244]^and_result1[245]^and_result1[246]^and_result1[247]^and_result1[248]^and_result1[249]^and_result1[250]^and_result1[251]^and_result1[252]^and_result1[253]^and_result1[254];
assign key[2]=and_result2[0]^and_result2[1]^and_result2[2]^and_result2[3]^and_result2[4]^and_result2[5]^and_result2[6]^and_result2[7]^and_result2[8]^and_result2[9]^and_result2[10]^and_result2[11]^and_result2[12]^and_result2[13]^and_result2[14]^and_result2[15]^and_result2[16]^and_result2[17]^and_result2[18]^and_result2[19]^and_result2[20]^and_result2[21]^and_result2[22]^and_result2[23]^and_result2[24]^and_result2[25]^and_result2[26]^and_result2[27]^and_result2[28]^and_result2[29]^and_result2[30]^and_result2[31]^and_result2[32]^and_result2[33]^and_result2[34]^and_result2[35]^and_result2[36]^and_result2[37]^and_result2[38]^and_result2[39]^and_result2[40]^and_result2[41]^and_result2[42]^and_result2[43]^and_result2[44]^and_result2[45]^and_result2[46]^and_result2[47]^and_result2[48]^and_result2[49]^and_result2[50]^and_result2[51]^and_result2[52]^and_result2[53]^and_result2[54]^and_result2[55]^and_result2[56]^and_result2[57]^and_result2[58]^and_result2[59]^and_result2[60]^and_result2[61]^and_result2[62]^and_result2[63]^and_result2[64]^and_result2[65]^and_result2[66]^and_result2[67]^and_result2[68]^and_result2[69]^and_result2[70]^and_result2[71]^and_result2[72]^and_result2[73]^and_result2[74]^and_result2[75]^and_result2[76]^and_result2[77]^and_result2[78]^and_result2[79]^and_result2[80]^and_result2[81]^and_result2[82]^and_result2[83]^and_result2[84]^and_result2[85]^and_result2[86]^and_result2[87]^and_result2[88]^and_result2[89]^and_result2[90]^and_result2[91]^and_result2[92]^and_result2[93]^and_result2[94]^and_result2[95]^and_result2[96]^and_result2[97]^and_result2[98]^and_result2[99]^and_result2[100]^and_result2[101]^and_result2[102]^and_result2[103]^and_result2[104]^and_result2[105]^and_result2[106]^and_result2[107]^and_result2[108]^and_result2[109]^and_result2[110]^and_result2[111]^and_result2[112]^and_result2[113]^and_result2[114]^and_result2[115]^and_result2[116]^and_result2[117]^and_result2[118]^and_result2[119]^and_result2[120]^and_result2[121]^and_result2[122]^and_result2[123]^and_result2[124]^and_result2[125]^and_result2[126]^and_result2[127]^and_result2[128]^and_result2[129]^and_result2[130]^and_result2[131]^and_result2[132]^and_result2[133]^and_result2[134]^and_result2[135]^and_result2[136]^and_result2[137]^and_result2[138]^and_result2[139]^and_result2[140]^and_result2[141]^and_result2[142]^and_result2[143]^and_result2[144]^and_result2[145]^and_result2[146]^and_result2[147]^and_result2[148]^and_result2[149]^and_result2[150]^and_result2[151]^and_result2[152]^and_result2[153]^and_result2[154]^and_result2[155]^and_result2[156]^and_result2[157]^and_result2[158]^and_result2[159]^and_result2[160]^and_result2[161]^and_result2[162]^and_result2[163]^and_result2[164]^and_result2[165]^and_result2[166]^and_result2[167]^and_result2[168]^and_result2[169]^and_result2[170]^and_result2[171]^and_result2[172]^and_result2[173]^and_result2[174]^and_result2[175]^and_result2[176]^and_result2[177]^and_result2[178]^and_result2[179]^and_result2[180]^and_result2[181]^and_result2[182]^and_result2[183]^and_result2[184]^and_result2[185]^and_result2[186]^and_result2[187]^and_result2[188]^and_result2[189]^and_result2[190]^and_result2[191]^and_result2[192]^and_result2[193]^and_result2[194]^and_result2[195]^and_result2[196]^and_result2[197]^and_result2[198]^and_result2[199]^and_result2[200]^and_result2[201]^and_result2[202]^and_result2[203]^and_result2[204]^and_result2[205]^and_result2[206]^and_result2[207]^and_result2[208]^and_result2[209]^and_result2[210]^and_result2[211]^and_result2[212]^and_result2[213]^and_result2[214]^and_result2[215]^and_result2[216]^and_result2[217]^and_result2[218]^and_result2[219]^and_result2[220]^and_result2[221]^and_result2[222]^and_result2[223]^and_result2[224]^and_result2[225]^and_result2[226]^and_result2[227]^and_result2[228]^and_result2[229]^and_result2[230]^and_result2[231]^and_result2[232]^and_result2[233]^and_result2[234]^and_result2[235]^and_result2[236]^and_result2[237]^and_result2[238]^and_result2[239]^and_result2[240]^and_result2[241]^and_result2[242]^and_result2[243]^and_result2[244]^and_result2[245]^and_result2[246]^and_result2[247]^and_result2[248]^and_result2[249]^and_result2[250]^and_result2[251]^and_result2[252]^and_result2[253]^and_result2[254];
assign key[3]=and_result3[0]^and_result3[1]^and_result3[2]^and_result3[3]^and_result3[4]^and_result3[5]^and_result3[6]^and_result3[7]^and_result3[8]^and_result3[9]^and_result3[10]^and_result3[11]^and_result3[12]^and_result3[13]^and_result3[14]^and_result3[15]^and_result3[16]^and_result3[17]^and_result3[18]^and_result3[19]^and_result3[20]^and_result3[21]^and_result3[22]^and_result3[23]^and_result3[24]^and_result3[25]^and_result3[26]^and_result3[27]^and_result3[28]^and_result3[29]^and_result3[30]^and_result3[31]^and_result3[32]^and_result3[33]^and_result3[34]^and_result3[35]^and_result3[36]^and_result3[37]^and_result3[38]^and_result3[39]^and_result3[40]^and_result3[41]^and_result3[42]^and_result3[43]^and_result3[44]^and_result3[45]^and_result3[46]^and_result3[47]^and_result3[48]^and_result3[49]^and_result3[50]^and_result3[51]^and_result3[52]^and_result3[53]^and_result3[54]^and_result3[55]^and_result3[56]^and_result3[57]^and_result3[58]^and_result3[59]^and_result3[60]^and_result3[61]^and_result3[62]^and_result3[63]^and_result3[64]^and_result3[65]^and_result3[66]^and_result3[67]^and_result3[68]^and_result3[69]^and_result3[70]^and_result3[71]^and_result3[72]^and_result3[73]^and_result3[74]^and_result3[75]^and_result3[76]^and_result3[77]^and_result3[78]^and_result3[79]^and_result3[80]^and_result3[81]^and_result3[82]^and_result3[83]^and_result3[84]^and_result3[85]^and_result3[86]^and_result3[87]^and_result3[88]^and_result3[89]^and_result3[90]^and_result3[91]^and_result3[92]^and_result3[93]^and_result3[94]^and_result3[95]^and_result3[96]^and_result3[97]^and_result3[98]^and_result3[99]^and_result3[100]^and_result3[101]^and_result3[102]^and_result3[103]^and_result3[104]^and_result3[105]^and_result3[106]^and_result3[107]^and_result3[108]^and_result3[109]^and_result3[110]^and_result3[111]^and_result3[112]^and_result3[113]^and_result3[114]^and_result3[115]^and_result3[116]^and_result3[117]^and_result3[118]^and_result3[119]^and_result3[120]^and_result3[121]^and_result3[122]^and_result3[123]^and_result3[124]^and_result3[125]^and_result3[126]^and_result3[127]^and_result3[128]^and_result3[129]^and_result3[130]^and_result3[131]^and_result3[132]^and_result3[133]^and_result3[134]^and_result3[135]^and_result3[136]^and_result3[137]^and_result3[138]^and_result3[139]^and_result3[140]^and_result3[141]^and_result3[142]^and_result3[143]^and_result3[144]^and_result3[145]^and_result3[146]^and_result3[147]^and_result3[148]^and_result3[149]^and_result3[150]^and_result3[151]^and_result3[152]^and_result3[153]^and_result3[154]^and_result3[155]^and_result3[156]^and_result3[157]^and_result3[158]^and_result3[159]^and_result3[160]^and_result3[161]^and_result3[162]^and_result3[163]^and_result3[164]^and_result3[165]^and_result3[166]^and_result3[167]^and_result3[168]^and_result3[169]^and_result3[170]^and_result3[171]^and_result3[172]^and_result3[173]^and_result3[174]^and_result3[175]^and_result3[176]^and_result3[177]^and_result3[178]^and_result3[179]^and_result3[180]^and_result3[181]^and_result3[182]^and_result3[183]^and_result3[184]^and_result3[185]^and_result3[186]^and_result3[187]^and_result3[188]^and_result3[189]^and_result3[190]^and_result3[191]^and_result3[192]^and_result3[193]^and_result3[194]^and_result3[195]^and_result3[196]^and_result3[197]^and_result3[198]^and_result3[199]^and_result3[200]^and_result3[201]^and_result3[202]^and_result3[203]^and_result3[204]^and_result3[205]^and_result3[206]^and_result3[207]^and_result3[208]^and_result3[209]^and_result3[210]^and_result3[211]^and_result3[212]^and_result3[213]^and_result3[214]^and_result3[215]^and_result3[216]^and_result3[217]^and_result3[218]^and_result3[219]^and_result3[220]^and_result3[221]^and_result3[222]^and_result3[223]^and_result3[224]^and_result3[225]^and_result3[226]^and_result3[227]^and_result3[228]^and_result3[229]^and_result3[230]^and_result3[231]^and_result3[232]^and_result3[233]^and_result3[234]^and_result3[235]^and_result3[236]^and_result3[237]^and_result3[238]^and_result3[239]^and_result3[240]^and_result3[241]^and_result3[242]^and_result3[243]^and_result3[244]^and_result3[245]^and_result3[246]^and_result3[247]^and_result3[248]^and_result3[249]^and_result3[250]^and_result3[251]^and_result3[252]^and_result3[253]^and_result3[254];
assign key[4]=and_result4[0]^and_result4[1]^and_result4[2]^and_result4[3]^and_result4[4]^and_result4[5]^and_result4[6]^and_result4[7]^and_result4[8]^and_result4[9]^and_result4[10]^and_result4[11]^and_result4[12]^and_result4[13]^and_result4[14]^and_result4[15]^and_result4[16]^and_result4[17]^and_result4[18]^and_result4[19]^and_result4[20]^and_result4[21]^and_result4[22]^and_result4[23]^and_result4[24]^and_result4[25]^and_result4[26]^and_result4[27]^and_result4[28]^and_result4[29]^and_result4[30]^and_result4[31]^and_result4[32]^and_result4[33]^and_result4[34]^and_result4[35]^and_result4[36]^and_result4[37]^and_result4[38]^and_result4[39]^and_result4[40]^and_result4[41]^and_result4[42]^and_result4[43]^and_result4[44]^and_result4[45]^and_result4[46]^and_result4[47]^and_result4[48]^and_result4[49]^and_result4[50]^and_result4[51]^and_result4[52]^and_result4[53]^and_result4[54]^and_result4[55]^and_result4[56]^and_result4[57]^and_result4[58]^and_result4[59]^and_result4[60]^and_result4[61]^and_result4[62]^and_result4[63]^and_result4[64]^and_result4[65]^and_result4[66]^and_result4[67]^and_result4[68]^and_result4[69]^and_result4[70]^and_result4[71]^and_result4[72]^and_result4[73]^and_result4[74]^and_result4[75]^and_result4[76]^and_result4[77]^and_result4[78]^and_result4[79]^and_result4[80]^and_result4[81]^and_result4[82]^and_result4[83]^and_result4[84]^and_result4[85]^and_result4[86]^and_result4[87]^and_result4[88]^and_result4[89]^and_result4[90]^and_result4[91]^and_result4[92]^and_result4[93]^and_result4[94]^and_result4[95]^and_result4[96]^and_result4[97]^and_result4[98]^and_result4[99]^and_result4[100]^and_result4[101]^and_result4[102]^and_result4[103]^and_result4[104]^and_result4[105]^and_result4[106]^and_result4[107]^and_result4[108]^and_result4[109]^and_result4[110]^and_result4[111]^and_result4[112]^and_result4[113]^and_result4[114]^and_result4[115]^and_result4[116]^and_result4[117]^and_result4[118]^and_result4[119]^and_result4[120]^and_result4[121]^and_result4[122]^and_result4[123]^and_result4[124]^and_result4[125]^and_result4[126]^and_result4[127]^and_result4[128]^and_result4[129]^and_result4[130]^and_result4[131]^and_result4[132]^and_result4[133]^and_result4[134]^and_result4[135]^and_result4[136]^and_result4[137]^and_result4[138]^and_result4[139]^and_result4[140]^and_result4[141]^and_result4[142]^and_result4[143]^and_result4[144]^and_result4[145]^and_result4[146]^and_result4[147]^and_result4[148]^and_result4[149]^and_result4[150]^and_result4[151]^and_result4[152]^and_result4[153]^and_result4[154]^and_result4[155]^and_result4[156]^and_result4[157]^and_result4[158]^and_result4[159]^and_result4[160]^and_result4[161]^and_result4[162]^and_result4[163]^and_result4[164]^and_result4[165]^and_result4[166]^and_result4[167]^and_result4[168]^and_result4[169]^and_result4[170]^and_result4[171]^and_result4[172]^and_result4[173]^and_result4[174]^and_result4[175]^and_result4[176]^and_result4[177]^and_result4[178]^and_result4[179]^and_result4[180]^and_result4[181]^and_result4[182]^and_result4[183]^and_result4[184]^and_result4[185]^and_result4[186]^and_result4[187]^and_result4[188]^and_result4[189]^and_result4[190]^and_result4[191]^and_result4[192]^and_result4[193]^and_result4[194]^and_result4[195]^and_result4[196]^and_result4[197]^and_result4[198]^and_result4[199]^and_result4[200]^and_result4[201]^and_result4[202]^and_result4[203]^and_result4[204]^and_result4[205]^and_result4[206]^and_result4[207]^and_result4[208]^and_result4[209]^and_result4[210]^and_result4[211]^and_result4[212]^and_result4[213]^and_result4[214]^and_result4[215]^and_result4[216]^and_result4[217]^and_result4[218]^and_result4[219]^and_result4[220]^and_result4[221]^and_result4[222]^and_result4[223]^and_result4[224]^and_result4[225]^and_result4[226]^and_result4[227]^and_result4[228]^and_result4[229]^and_result4[230]^and_result4[231]^and_result4[232]^and_result4[233]^and_result4[234]^and_result4[235]^and_result4[236]^and_result4[237]^and_result4[238]^and_result4[239]^and_result4[240]^and_result4[241]^and_result4[242]^and_result4[243]^and_result4[244]^and_result4[245]^and_result4[246]^and_result4[247]^and_result4[248]^and_result4[249]^and_result4[250]^and_result4[251]^and_result4[252]^and_result4[253]^and_result4[254];
assign key[5]=and_result5[0]^and_result5[1]^and_result5[2]^and_result5[3]^and_result5[4]^and_result5[5]^and_result5[6]^and_result5[7]^and_result5[8]^and_result5[9]^and_result5[10]^and_result5[11]^and_result5[12]^and_result5[13]^and_result5[14]^and_result5[15]^and_result5[16]^and_result5[17]^and_result5[18]^and_result5[19]^and_result5[20]^and_result5[21]^and_result5[22]^and_result5[23]^and_result5[24]^and_result5[25]^and_result5[26]^and_result5[27]^and_result5[28]^and_result5[29]^and_result5[30]^and_result5[31]^and_result5[32]^and_result5[33]^and_result5[34]^and_result5[35]^and_result5[36]^and_result5[37]^and_result5[38]^and_result5[39]^and_result5[40]^and_result5[41]^and_result5[42]^and_result5[43]^and_result5[44]^and_result5[45]^and_result5[46]^and_result5[47]^and_result5[48]^and_result5[49]^and_result5[50]^and_result5[51]^and_result5[52]^and_result5[53]^and_result5[54]^and_result5[55]^and_result5[56]^and_result5[57]^and_result5[58]^and_result5[59]^and_result5[60]^and_result5[61]^and_result5[62]^and_result5[63]^and_result5[64]^and_result5[65]^and_result5[66]^and_result5[67]^and_result5[68]^and_result5[69]^and_result5[70]^and_result5[71]^and_result5[72]^and_result5[73]^and_result5[74]^and_result5[75]^and_result5[76]^and_result5[77]^and_result5[78]^and_result5[79]^and_result5[80]^and_result5[81]^and_result5[82]^and_result5[83]^and_result5[84]^and_result5[85]^and_result5[86]^and_result5[87]^and_result5[88]^and_result5[89]^and_result5[90]^and_result5[91]^and_result5[92]^and_result5[93]^and_result5[94]^and_result5[95]^and_result5[96]^and_result5[97]^and_result5[98]^and_result5[99]^and_result5[100]^and_result5[101]^and_result5[102]^and_result5[103]^and_result5[104]^and_result5[105]^and_result5[106]^and_result5[107]^and_result5[108]^and_result5[109]^and_result5[110]^and_result5[111]^and_result5[112]^and_result5[113]^and_result5[114]^and_result5[115]^and_result5[116]^and_result5[117]^and_result5[118]^and_result5[119]^and_result5[120]^and_result5[121]^and_result5[122]^and_result5[123]^and_result5[124]^and_result5[125]^and_result5[126]^and_result5[127]^and_result5[128]^and_result5[129]^and_result5[130]^and_result5[131]^and_result5[132]^and_result5[133]^and_result5[134]^and_result5[135]^and_result5[136]^and_result5[137]^and_result5[138]^and_result5[139]^and_result5[140]^and_result5[141]^and_result5[142]^and_result5[143]^and_result5[144]^and_result5[145]^and_result5[146]^and_result5[147]^and_result5[148]^and_result5[149]^and_result5[150]^and_result5[151]^and_result5[152]^and_result5[153]^and_result5[154]^and_result5[155]^and_result5[156]^and_result5[157]^and_result5[158]^and_result5[159]^and_result5[160]^and_result5[161]^and_result5[162]^and_result5[163]^and_result5[164]^and_result5[165]^and_result5[166]^and_result5[167]^and_result5[168]^and_result5[169]^and_result5[170]^and_result5[171]^and_result5[172]^and_result5[173]^and_result5[174]^and_result5[175]^and_result5[176]^and_result5[177]^and_result5[178]^and_result5[179]^and_result5[180]^and_result5[181]^and_result5[182]^and_result5[183]^and_result5[184]^and_result5[185]^and_result5[186]^and_result5[187]^and_result5[188]^and_result5[189]^and_result5[190]^and_result5[191]^and_result5[192]^and_result5[193]^and_result5[194]^and_result5[195]^and_result5[196]^and_result5[197]^and_result5[198]^and_result5[199]^and_result5[200]^and_result5[201]^and_result5[202]^and_result5[203]^and_result5[204]^and_result5[205]^and_result5[206]^and_result5[207]^and_result5[208]^and_result5[209]^and_result5[210]^and_result5[211]^and_result5[212]^and_result5[213]^and_result5[214]^and_result5[215]^and_result5[216]^and_result5[217]^and_result5[218]^and_result5[219]^and_result5[220]^and_result5[221]^and_result5[222]^and_result5[223]^and_result5[224]^and_result5[225]^and_result5[226]^and_result5[227]^and_result5[228]^and_result5[229]^and_result5[230]^and_result5[231]^and_result5[232]^and_result5[233]^and_result5[234]^and_result5[235]^and_result5[236]^and_result5[237]^and_result5[238]^and_result5[239]^and_result5[240]^and_result5[241]^and_result5[242]^and_result5[243]^and_result5[244]^and_result5[245]^and_result5[246]^and_result5[247]^and_result5[248]^and_result5[249]^and_result5[250]^and_result5[251]^and_result5[252]^and_result5[253]^and_result5[254];
assign key[6]=and_result6[0]^and_result6[1]^and_result6[2]^and_result6[3]^and_result6[4]^and_result6[5]^and_result6[6]^and_result6[7]^and_result6[8]^and_result6[9]^and_result6[10]^and_result6[11]^and_result6[12]^and_result6[13]^and_result6[14]^and_result6[15]^and_result6[16]^and_result6[17]^and_result6[18]^and_result6[19]^and_result6[20]^and_result6[21]^and_result6[22]^and_result6[23]^and_result6[24]^and_result6[25]^and_result6[26]^and_result6[27]^and_result6[28]^and_result6[29]^and_result6[30]^and_result6[31]^and_result6[32]^and_result6[33]^and_result6[34]^and_result6[35]^and_result6[36]^and_result6[37]^and_result6[38]^and_result6[39]^and_result6[40]^and_result6[41]^and_result6[42]^and_result6[43]^and_result6[44]^and_result6[45]^and_result6[46]^and_result6[47]^and_result6[48]^and_result6[49]^and_result6[50]^and_result6[51]^and_result6[52]^and_result6[53]^and_result6[54]^and_result6[55]^and_result6[56]^and_result6[57]^and_result6[58]^and_result6[59]^and_result6[60]^and_result6[61]^and_result6[62]^and_result6[63]^and_result6[64]^and_result6[65]^and_result6[66]^and_result6[67]^and_result6[68]^and_result6[69]^and_result6[70]^and_result6[71]^and_result6[72]^and_result6[73]^and_result6[74]^and_result6[75]^and_result6[76]^and_result6[77]^and_result6[78]^and_result6[79]^and_result6[80]^and_result6[81]^and_result6[82]^and_result6[83]^and_result6[84]^and_result6[85]^and_result6[86]^and_result6[87]^and_result6[88]^and_result6[89]^and_result6[90]^and_result6[91]^and_result6[92]^and_result6[93]^and_result6[94]^and_result6[95]^and_result6[96]^and_result6[97]^and_result6[98]^and_result6[99]^and_result6[100]^and_result6[101]^and_result6[102]^and_result6[103]^and_result6[104]^and_result6[105]^and_result6[106]^and_result6[107]^and_result6[108]^and_result6[109]^and_result6[110]^and_result6[111]^and_result6[112]^and_result6[113]^and_result6[114]^and_result6[115]^and_result6[116]^and_result6[117]^and_result6[118]^and_result6[119]^and_result6[120]^and_result6[121]^and_result6[122]^and_result6[123]^and_result6[124]^and_result6[125]^and_result6[126]^and_result6[127]^and_result6[128]^and_result6[129]^and_result6[130]^and_result6[131]^and_result6[132]^and_result6[133]^and_result6[134]^and_result6[135]^and_result6[136]^and_result6[137]^and_result6[138]^and_result6[139]^and_result6[140]^and_result6[141]^and_result6[142]^and_result6[143]^and_result6[144]^and_result6[145]^and_result6[146]^and_result6[147]^and_result6[148]^and_result6[149]^and_result6[150]^and_result6[151]^and_result6[152]^and_result6[153]^and_result6[154]^and_result6[155]^and_result6[156]^and_result6[157]^and_result6[158]^and_result6[159]^and_result6[160]^and_result6[161]^and_result6[162]^and_result6[163]^and_result6[164]^and_result6[165]^and_result6[166]^and_result6[167]^and_result6[168]^and_result6[169]^and_result6[170]^and_result6[171]^and_result6[172]^and_result6[173]^and_result6[174]^and_result6[175]^and_result6[176]^and_result6[177]^and_result6[178]^and_result6[179]^and_result6[180]^and_result6[181]^and_result6[182]^and_result6[183]^and_result6[184]^and_result6[185]^and_result6[186]^and_result6[187]^and_result6[188]^and_result6[189]^and_result6[190]^and_result6[191]^and_result6[192]^and_result6[193]^and_result6[194]^and_result6[195]^and_result6[196]^and_result6[197]^and_result6[198]^and_result6[199]^and_result6[200]^and_result6[201]^and_result6[202]^and_result6[203]^and_result6[204]^and_result6[205]^and_result6[206]^and_result6[207]^and_result6[208]^and_result6[209]^and_result6[210]^and_result6[211]^and_result6[212]^and_result6[213]^and_result6[214]^and_result6[215]^and_result6[216]^and_result6[217]^and_result6[218]^and_result6[219]^and_result6[220]^and_result6[221]^and_result6[222]^and_result6[223]^and_result6[224]^and_result6[225]^and_result6[226]^and_result6[227]^and_result6[228]^and_result6[229]^and_result6[230]^and_result6[231]^and_result6[232]^and_result6[233]^and_result6[234]^and_result6[235]^and_result6[236]^and_result6[237]^and_result6[238]^and_result6[239]^and_result6[240]^and_result6[241]^and_result6[242]^and_result6[243]^and_result6[244]^and_result6[245]^and_result6[246]^and_result6[247]^and_result6[248]^and_result6[249]^and_result6[250]^and_result6[251]^and_result6[252]^and_result6[253]^and_result6[254];
assign key[7]=and_result7[0]^and_result7[1]^and_result7[2]^and_result7[3]^and_result7[4]^and_result7[5]^and_result7[6]^and_result7[7]^and_result7[8]^and_result7[9]^and_result7[10]^and_result7[11]^and_result7[12]^and_result7[13]^and_result7[14]^and_result7[15]^and_result7[16]^and_result7[17]^and_result7[18]^and_result7[19]^and_result7[20]^and_result7[21]^and_result7[22]^and_result7[23]^and_result7[24]^and_result7[25]^and_result7[26]^and_result7[27]^and_result7[28]^and_result7[29]^and_result7[30]^and_result7[31]^and_result7[32]^and_result7[33]^and_result7[34]^and_result7[35]^and_result7[36]^and_result7[37]^and_result7[38]^and_result7[39]^and_result7[40]^and_result7[41]^and_result7[42]^and_result7[43]^and_result7[44]^and_result7[45]^and_result7[46]^and_result7[47]^and_result7[48]^and_result7[49]^and_result7[50]^and_result7[51]^and_result7[52]^and_result7[53]^and_result7[54]^and_result7[55]^and_result7[56]^and_result7[57]^and_result7[58]^and_result7[59]^and_result7[60]^and_result7[61]^and_result7[62]^and_result7[63]^and_result7[64]^and_result7[65]^and_result7[66]^and_result7[67]^and_result7[68]^and_result7[69]^and_result7[70]^and_result7[71]^and_result7[72]^and_result7[73]^and_result7[74]^and_result7[75]^and_result7[76]^and_result7[77]^and_result7[78]^and_result7[79]^and_result7[80]^and_result7[81]^and_result7[82]^and_result7[83]^and_result7[84]^and_result7[85]^and_result7[86]^and_result7[87]^and_result7[88]^and_result7[89]^and_result7[90]^and_result7[91]^and_result7[92]^and_result7[93]^and_result7[94]^and_result7[95]^and_result7[96]^and_result7[97]^and_result7[98]^and_result7[99]^and_result7[100]^and_result7[101]^and_result7[102]^and_result7[103]^and_result7[104]^and_result7[105]^and_result7[106]^and_result7[107]^and_result7[108]^and_result7[109]^and_result7[110]^and_result7[111]^and_result7[112]^and_result7[113]^and_result7[114]^and_result7[115]^and_result7[116]^and_result7[117]^and_result7[118]^and_result7[119]^and_result7[120]^and_result7[121]^and_result7[122]^and_result7[123]^and_result7[124]^and_result7[125]^and_result7[126]^and_result7[127]^and_result7[128]^and_result7[129]^and_result7[130]^and_result7[131]^and_result7[132]^and_result7[133]^and_result7[134]^and_result7[135]^and_result7[136]^and_result7[137]^and_result7[138]^and_result7[139]^and_result7[140]^and_result7[141]^and_result7[142]^and_result7[143]^and_result7[144]^and_result7[145]^and_result7[146]^and_result7[147]^and_result7[148]^and_result7[149]^and_result7[150]^and_result7[151]^and_result7[152]^and_result7[153]^and_result7[154]^and_result7[155]^and_result7[156]^and_result7[157]^and_result7[158]^and_result7[159]^and_result7[160]^and_result7[161]^and_result7[162]^and_result7[163]^and_result7[164]^and_result7[165]^and_result7[166]^and_result7[167]^and_result7[168]^and_result7[169]^and_result7[170]^and_result7[171]^and_result7[172]^and_result7[173]^and_result7[174]^and_result7[175]^and_result7[176]^and_result7[177]^and_result7[178]^and_result7[179]^and_result7[180]^and_result7[181]^and_result7[182]^and_result7[183]^and_result7[184]^and_result7[185]^and_result7[186]^and_result7[187]^and_result7[188]^and_result7[189]^and_result7[190]^and_result7[191]^and_result7[192]^and_result7[193]^and_result7[194]^and_result7[195]^and_result7[196]^and_result7[197]^and_result7[198]^and_result7[199]^and_result7[200]^and_result7[201]^and_result7[202]^and_result7[203]^and_result7[204]^and_result7[205]^and_result7[206]^and_result7[207]^and_result7[208]^and_result7[209]^and_result7[210]^and_result7[211]^and_result7[212]^and_result7[213]^and_result7[214]^and_result7[215]^and_result7[216]^and_result7[217]^and_result7[218]^and_result7[219]^and_result7[220]^and_result7[221]^and_result7[222]^and_result7[223]^and_result7[224]^and_result7[225]^and_result7[226]^and_result7[227]^and_result7[228]^and_result7[229]^and_result7[230]^and_result7[231]^and_result7[232]^and_result7[233]^and_result7[234]^and_result7[235]^and_result7[236]^and_result7[237]^and_result7[238]^and_result7[239]^and_result7[240]^and_result7[241]^and_result7[242]^and_result7[243]^and_result7[244]^and_result7[245]^and_result7[246]^and_result7[247]^and_result7[248]^and_result7[249]^and_result7[250]^and_result7[251]^and_result7[252]^and_result7[253]^and_result7[254];
assign key[8]=and_result8[0]^and_result8[1]^and_result8[2]^and_result8[3]^and_result8[4]^and_result8[5]^and_result8[6]^and_result8[7]^and_result8[8]^and_result8[9]^and_result8[10]^and_result8[11]^and_result8[12]^and_result8[13]^and_result8[14]^and_result8[15]^and_result8[16]^and_result8[17]^and_result8[18]^and_result8[19]^and_result8[20]^and_result8[21]^and_result8[22]^and_result8[23]^and_result8[24]^and_result8[25]^and_result8[26]^and_result8[27]^and_result8[28]^and_result8[29]^and_result8[30]^and_result8[31]^and_result8[32]^and_result8[33]^and_result8[34]^and_result8[35]^and_result8[36]^and_result8[37]^and_result8[38]^and_result8[39]^and_result8[40]^and_result8[41]^and_result8[42]^and_result8[43]^and_result8[44]^and_result8[45]^and_result8[46]^and_result8[47]^and_result8[48]^and_result8[49]^and_result8[50]^and_result8[51]^and_result8[52]^and_result8[53]^and_result8[54]^and_result8[55]^and_result8[56]^and_result8[57]^and_result8[58]^and_result8[59]^and_result8[60]^and_result8[61]^and_result8[62]^and_result8[63]^and_result8[64]^and_result8[65]^and_result8[66]^and_result8[67]^and_result8[68]^and_result8[69]^and_result8[70]^and_result8[71]^and_result8[72]^and_result8[73]^and_result8[74]^and_result8[75]^and_result8[76]^and_result8[77]^and_result8[78]^and_result8[79]^and_result8[80]^and_result8[81]^and_result8[82]^and_result8[83]^and_result8[84]^and_result8[85]^and_result8[86]^and_result8[87]^and_result8[88]^and_result8[89]^and_result8[90]^and_result8[91]^and_result8[92]^and_result8[93]^and_result8[94]^and_result8[95]^and_result8[96]^and_result8[97]^and_result8[98]^and_result8[99]^and_result8[100]^and_result8[101]^and_result8[102]^and_result8[103]^and_result8[104]^and_result8[105]^and_result8[106]^and_result8[107]^and_result8[108]^and_result8[109]^and_result8[110]^and_result8[111]^and_result8[112]^and_result8[113]^and_result8[114]^and_result8[115]^and_result8[116]^and_result8[117]^and_result8[118]^and_result8[119]^and_result8[120]^and_result8[121]^and_result8[122]^and_result8[123]^and_result8[124]^and_result8[125]^and_result8[126]^and_result8[127]^and_result8[128]^and_result8[129]^and_result8[130]^and_result8[131]^and_result8[132]^and_result8[133]^and_result8[134]^and_result8[135]^and_result8[136]^and_result8[137]^and_result8[138]^and_result8[139]^and_result8[140]^and_result8[141]^and_result8[142]^and_result8[143]^and_result8[144]^and_result8[145]^and_result8[146]^and_result8[147]^and_result8[148]^and_result8[149]^and_result8[150]^and_result8[151]^and_result8[152]^and_result8[153]^and_result8[154]^and_result8[155]^and_result8[156]^and_result8[157]^and_result8[158]^and_result8[159]^and_result8[160]^and_result8[161]^and_result8[162]^and_result8[163]^and_result8[164]^and_result8[165]^and_result8[166]^and_result8[167]^and_result8[168]^and_result8[169]^and_result8[170]^and_result8[171]^and_result8[172]^and_result8[173]^and_result8[174]^and_result8[175]^and_result8[176]^and_result8[177]^and_result8[178]^and_result8[179]^and_result8[180]^and_result8[181]^and_result8[182]^and_result8[183]^and_result8[184]^and_result8[185]^and_result8[186]^and_result8[187]^and_result8[188]^and_result8[189]^and_result8[190]^and_result8[191]^and_result8[192]^and_result8[193]^and_result8[194]^and_result8[195]^and_result8[196]^and_result8[197]^and_result8[198]^and_result8[199]^and_result8[200]^and_result8[201]^and_result8[202]^and_result8[203]^and_result8[204]^and_result8[205]^and_result8[206]^and_result8[207]^and_result8[208]^and_result8[209]^and_result8[210]^and_result8[211]^and_result8[212]^and_result8[213]^and_result8[214]^and_result8[215]^and_result8[216]^and_result8[217]^and_result8[218]^and_result8[219]^and_result8[220]^and_result8[221]^and_result8[222]^and_result8[223]^and_result8[224]^and_result8[225]^and_result8[226]^and_result8[227]^and_result8[228]^and_result8[229]^and_result8[230]^and_result8[231]^and_result8[232]^and_result8[233]^and_result8[234]^and_result8[235]^and_result8[236]^and_result8[237]^and_result8[238]^and_result8[239]^and_result8[240]^and_result8[241]^and_result8[242]^and_result8[243]^and_result8[244]^and_result8[245]^and_result8[246]^and_result8[247]^and_result8[248]^and_result8[249]^and_result8[250]^and_result8[251]^and_result8[252]^and_result8[253]^and_result8[254];
assign key[9]=and_result9[0]^and_result9[1]^and_result9[2]^and_result9[3]^and_result9[4]^and_result9[5]^and_result9[6]^and_result9[7]^and_result9[8]^and_result9[9]^and_result9[10]^and_result9[11]^and_result9[12]^and_result9[13]^and_result9[14]^and_result9[15]^and_result9[16]^and_result9[17]^and_result9[18]^and_result9[19]^and_result9[20]^and_result9[21]^and_result9[22]^and_result9[23]^and_result9[24]^and_result9[25]^and_result9[26]^and_result9[27]^and_result9[28]^and_result9[29]^and_result9[30]^and_result9[31]^and_result9[32]^and_result9[33]^and_result9[34]^and_result9[35]^and_result9[36]^and_result9[37]^and_result9[38]^and_result9[39]^and_result9[40]^and_result9[41]^and_result9[42]^and_result9[43]^and_result9[44]^and_result9[45]^and_result9[46]^and_result9[47]^and_result9[48]^and_result9[49]^and_result9[50]^and_result9[51]^and_result9[52]^and_result9[53]^and_result9[54]^and_result9[55]^and_result9[56]^and_result9[57]^and_result9[58]^and_result9[59]^and_result9[60]^and_result9[61]^and_result9[62]^and_result9[63]^and_result9[64]^and_result9[65]^and_result9[66]^and_result9[67]^and_result9[68]^and_result9[69]^and_result9[70]^and_result9[71]^and_result9[72]^and_result9[73]^and_result9[74]^and_result9[75]^and_result9[76]^and_result9[77]^and_result9[78]^and_result9[79]^and_result9[80]^and_result9[81]^and_result9[82]^and_result9[83]^and_result9[84]^and_result9[85]^and_result9[86]^and_result9[87]^and_result9[88]^and_result9[89]^and_result9[90]^and_result9[91]^and_result9[92]^and_result9[93]^and_result9[94]^and_result9[95]^and_result9[96]^and_result9[97]^and_result9[98]^and_result9[99]^and_result9[100]^and_result9[101]^and_result9[102]^and_result9[103]^and_result9[104]^and_result9[105]^and_result9[106]^and_result9[107]^and_result9[108]^and_result9[109]^and_result9[110]^and_result9[111]^and_result9[112]^and_result9[113]^and_result9[114]^and_result9[115]^and_result9[116]^and_result9[117]^and_result9[118]^and_result9[119]^and_result9[120]^and_result9[121]^and_result9[122]^and_result9[123]^and_result9[124]^and_result9[125]^and_result9[126]^and_result9[127]^and_result9[128]^and_result9[129]^and_result9[130]^and_result9[131]^and_result9[132]^and_result9[133]^and_result9[134]^and_result9[135]^and_result9[136]^and_result9[137]^and_result9[138]^and_result9[139]^and_result9[140]^and_result9[141]^and_result9[142]^and_result9[143]^and_result9[144]^and_result9[145]^and_result9[146]^and_result9[147]^and_result9[148]^and_result9[149]^and_result9[150]^and_result9[151]^and_result9[152]^and_result9[153]^and_result9[154]^and_result9[155]^and_result9[156]^and_result9[157]^and_result9[158]^and_result9[159]^and_result9[160]^and_result9[161]^and_result9[162]^and_result9[163]^and_result9[164]^and_result9[165]^and_result9[166]^and_result9[167]^and_result9[168]^and_result9[169]^and_result9[170]^and_result9[171]^and_result9[172]^and_result9[173]^and_result9[174]^and_result9[175]^and_result9[176]^and_result9[177]^and_result9[178]^and_result9[179]^and_result9[180]^and_result9[181]^and_result9[182]^and_result9[183]^and_result9[184]^and_result9[185]^and_result9[186]^and_result9[187]^and_result9[188]^and_result9[189]^and_result9[190]^and_result9[191]^and_result9[192]^and_result9[193]^and_result9[194]^and_result9[195]^and_result9[196]^and_result9[197]^and_result9[198]^and_result9[199]^and_result9[200]^and_result9[201]^and_result9[202]^and_result9[203]^and_result9[204]^and_result9[205]^and_result9[206]^and_result9[207]^and_result9[208]^and_result9[209]^and_result9[210]^and_result9[211]^and_result9[212]^and_result9[213]^and_result9[214]^and_result9[215]^and_result9[216]^and_result9[217]^and_result9[218]^and_result9[219]^and_result9[220]^and_result9[221]^and_result9[222]^and_result9[223]^and_result9[224]^and_result9[225]^and_result9[226]^and_result9[227]^and_result9[228]^and_result9[229]^and_result9[230]^and_result9[231]^and_result9[232]^and_result9[233]^and_result9[234]^and_result9[235]^and_result9[236]^and_result9[237]^and_result9[238]^and_result9[239]^and_result9[240]^and_result9[241]^and_result9[242]^and_result9[243]^and_result9[244]^and_result9[245]^and_result9[246]^and_result9[247]^and_result9[248]^and_result9[249]^and_result9[250]^and_result9[251]^and_result9[252]^and_result9[253]^and_result9[254];
assign key[10]=and_result10[0]^and_result10[1]^and_result10[2]^and_result10[3]^and_result10[4]^and_result10[5]^and_result10[6]^and_result10[7]^and_result10[8]^and_result10[9]^and_result10[10]^and_result10[11]^and_result10[12]^and_result10[13]^and_result10[14]^and_result10[15]^and_result10[16]^and_result10[17]^and_result10[18]^and_result10[19]^and_result10[20]^and_result10[21]^and_result10[22]^and_result10[23]^and_result10[24]^and_result10[25]^and_result10[26]^and_result10[27]^and_result10[28]^and_result10[29]^and_result10[30]^and_result10[31]^and_result10[32]^and_result10[33]^and_result10[34]^and_result10[35]^and_result10[36]^and_result10[37]^and_result10[38]^and_result10[39]^and_result10[40]^and_result10[41]^and_result10[42]^and_result10[43]^and_result10[44]^and_result10[45]^and_result10[46]^and_result10[47]^and_result10[48]^and_result10[49]^and_result10[50]^and_result10[51]^and_result10[52]^and_result10[53]^and_result10[54]^and_result10[55]^and_result10[56]^and_result10[57]^and_result10[58]^and_result10[59]^and_result10[60]^and_result10[61]^and_result10[62]^and_result10[63]^and_result10[64]^and_result10[65]^and_result10[66]^and_result10[67]^and_result10[68]^and_result10[69]^and_result10[70]^and_result10[71]^and_result10[72]^and_result10[73]^and_result10[74]^and_result10[75]^and_result10[76]^and_result10[77]^and_result10[78]^and_result10[79]^and_result10[80]^and_result10[81]^and_result10[82]^and_result10[83]^and_result10[84]^and_result10[85]^and_result10[86]^and_result10[87]^and_result10[88]^and_result10[89]^and_result10[90]^and_result10[91]^and_result10[92]^and_result10[93]^and_result10[94]^and_result10[95]^and_result10[96]^and_result10[97]^and_result10[98]^and_result10[99]^and_result10[100]^and_result10[101]^and_result10[102]^and_result10[103]^and_result10[104]^and_result10[105]^and_result10[106]^and_result10[107]^and_result10[108]^and_result10[109]^and_result10[110]^and_result10[111]^and_result10[112]^and_result10[113]^and_result10[114]^and_result10[115]^and_result10[116]^and_result10[117]^and_result10[118]^and_result10[119]^and_result10[120]^and_result10[121]^and_result10[122]^and_result10[123]^and_result10[124]^and_result10[125]^and_result10[126]^and_result10[127]^and_result10[128]^and_result10[129]^and_result10[130]^and_result10[131]^and_result10[132]^and_result10[133]^and_result10[134]^and_result10[135]^and_result10[136]^and_result10[137]^and_result10[138]^and_result10[139]^and_result10[140]^and_result10[141]^and_result10[142]^and_result10[143]^and_result10[144]^and_result10[145]^and_result10[146]^and_result10[147]^and_result10[148]^and_result10[149]^and_result10[150]^and_result10[151]^and_result10[152]^and_result10[153]^and_result10[154]^and_result10[155]^and_result10[156]^and_result10[157]^and_result10[158]^and_result10[159]^and_result10[160]^and_result10[161]^and_result10[162]^and_result10[163]^and_result10[164]^and_result10[165]^and_result10[166]^and_result10[167]^and_result10[168]^and_result10[169]^and_result10[170]^and_result10[171]^and_result10[172]^and_result10[173]^and_result10[174]^and_result10[175]^and_result10[176]^and_result10[177]^and_result10[178]^and_result10[179]^and_result10[180]^and_result10[181]^and_result10[182]^and_result10[183]^and_result10[184]^and_result10[185]^and_result10[186]^and_result10[187]^and_result10[188]^and_result10[189]^and_result10[190]^and_result10[191]^and_result10[192]^and_result10[193]^and_result10[194]^and_result10[195]^and_result10[196]^and_result10[197]^and_result10[198]^and_result10[199]^and_result10[200]^and_result10[201]^and_result10[202]^and_result10[203]^and_result10[204]^and_result10[205]^and_result10[206]^and_result10[207]^and_result10[208]^and_result10[209]^and_result10[210]^and_result10[211]^and_result10[212]^and_result10[213]^and_result10[214]^and_result10[215]^and_result10[216]^and_result10[217]^and_result10[218]^and_result10[219]^and_result10[220]^and_result10[221]^and_result10[222]^and_result10[223]^and_result10[224]^and_result10[225]^and_result10[226]^and_result10[227]^and_result10[228]^and_result10[229]^and_result10[230]^and_result10[231]^and_result10[232]^and_result10[233]^and_result10[234]^and_result10[235]^and_result10[236]^and_result10[237]^and_result10[238]^and_result10[239]^and_result10[240]^and_result10[241]^and_result10[242]^and_result10[243]^and_result10[244]^and_result10[245]^and_result10[246]^and_result10[247]^and_result10[248]^and_result10[249]^and_result10[250]^and_result10[251]^and_result10[252]^and_result10[253]^and_result10[254];
assign key[11]=and_result11[0]^and_result11[1]^and_result11[2]^and_result11[3]^and_result11[4]^and_result11[5]^and_result11[6]^and_result11[7]^and_result11[8]^and_result11[9]^and_result11[10]^and_result11[11]^and_result11[12]^and_result11[13]^and_result11[14]^and_result11[15]^and_result11[16]^and_result11[17]^and_result11[18]^and_result11[19]^and_result11[20]^and_result11[21]^and_result11[22]^and_result11[23]^and_result11[24]^and_result11[25]^and_result11[26]^and_result11[27]^and_result11[28]^and_result11[29]^and_result11[30]^and_result11[31]^and_result11[32]^and_result11[33]^and_result11[34]^and_result11[35]^and_result11[36]^and_result11[37]^and_result11[38]^and_result11[39]^and_result11[40]^and_result11[41]^and_result11[42]^and_result11[43]^and_result11[44]^and_result11[45]^and_result11[46]^and_result11[47]^and_result11[48]^and_result11[49]^and_result11[50]^and_result11[51]^and_result11[52]^and_result11[53]^and_result11[54]^and_result11[55]^and_result11[56]^and_result11[57]^and_result11[58]^and_result11[59]^and_result11[60]^and_result11[61]^and_result11[62]^and_result11[63]^and_result11[64]^and_result11[65]^and_result11[66]^and_result11[67]^and_result11[68]^and_result11[69]^and_result11[70]^and_result11[71]^and_result11[72]^and_result11[73]^and_result11[74]^and_result11[75]^and_result11[76]^and_result11[77]^and_result11[78]^and_result11[79]^and_result11[80]^and_result11[81]^and_result11[82]^and_result11[83]^and_result11[84]^and_result11[85]^and_result11[86]^and_result11[87]^and_result11[88]^and_result11[89]^and_result11[90]^and_result11[91]^and_result11[92]^and_result11[93]^and_result11[94]^and_result11[95]^and_result11[96]^and_result11[97]^and_result11[98]^and_result11[99]^and_result11[100]^and_result11[101]^and_result11[102]^and_result11[103]^and_result11[104]^and_result11[105]^and_result11[106]^and_result11[107]^and_result11[108]^and_result11[109]^and_result11[110]^and_result11[111]^and_result11[112]^and_result11[113]^and_result11[114]^and_result11[115]^and_result11[116]^and_result11[117]^and_result11[118]^and_result11[119]^and_result11[120]^and_result11[121]^and_result11[122]^and_result11[123]^and_result11[124]^and_result11[125]^and_result11[126]^and_result11[127]^and_result11[128]^and_result11[129]^and_result11[130]^and_result11[131]^and_result11[132]^and_result11[133]^and_result11[134]^and_result11[135]^and_result11[136]^and_result11[137]^and_result11[138]^and_result11[139]^and_result11[140]^and_result11[141]^and_result11[142]^and_result11[143]^and_result11[144]^and_result11[145]^and_result11[146]^and_result11[147]^and_result11[148]^and_result11[149]^and_result11[150]^and_result11[151]^and_result11[152]^and_result11[153]^and_result11[154]^and_result11[155]^and_result11[156]^and_result11[157]^and_result11[158]^and_result11[159]^and_result11[160]^and_result11[161]^and_result11[162]^and_result11[163]^and_result11[164]^and_result11[165]^and_result11[166]^and_result11[167]^and_result11[168]^and_result11[169]^and_result11[170]^and_result11[171]^and_result11[172]^and_result11[173]^and_result11[174]^and_result11[175]^and_result11[176]^and_result11[177]^and_result11[178]^and_result11[179]^and_result11[180]^and_result11[181]^and_result11[182]^and_result11[183]^and_result11[184]^and_result11[185]^and_result11[186]^and_result11[187]^and_result11[188]^and_result11[189]^and_result11[190]^and_result11[191]^and_result11[192]^and_result11[193]^and_result11[194]^and_result11[195]^and_result11[196]^and_result11[197]^and_result11[198]^and_result11[199]^and_result11[200]^and_result11[201]^and_result11[202]^and_result11[203]^and_result11[204]^and_result11[205]^and_result11[206]^and_result11[207]^and_result11[208]^and_result11[209]^and_result11[210]^and_result11[211]^and_result11[212]^and_result11[213]^and_result11[214]^and_result11[215]^and_result11[216]^and_result11[217]^and_result11[218]^and_result11[219]^and_result11[220]^and_result11[221]^and_result11[222]^and_result11[223]^and_result11[224]^and_result11[225]^and_result11[226]^and_result11[227]^and_result11[228]^and_result11[229]^and_result11[230]^and_result11[231]^and_result11[232]^and_result11[233]^and_result11[234]^and_result11[235]^and_result11[236]^and_result11[237]^and_result11[238]^and_result11[239]^and_result11[240]^and_result11[241]^and_result11[242]^and_result11[243]^and_result11[244]^and_result11[245]^and_result11[246]^and_result11[247]^and_result11[248]^and_result11[249]^and_result11[250]^and_result11[251]^and_result11[252]^and_result11[253]^and_result11[254];
assign key[12]=and_result12[0]^and_result12[1]^and_result12[2]^and_result12[3]^and_result12[4]^and_result12[5]^and_result12[6]^and_result12[7]^and_result12[8]^and_result12[9]^and_result12[10]^and_result12[11]^and_result12[12]^and_result12[13]^and_result12[14]^and_result12[15]^and_result12[16]^and_result12[17]^and_result12[18]^and_result12[19]^and_result12[20]^and_result12[21]^and_result12[22]^and_result12[23]^and_result12[24]^and_result12[25]^and_result12[26]^and_result12[27]^and_result12[28]^and_result12[29]^and_result12[30]^and_result12[31]^and_result12[32]^and_result12[33]^and_result12[34]^and_result12[35]^and_result12[36]^and_result12[37]^and_result12[38]^and_result12[39]^and_result12[40]^and_result12[41]^and_result12[42]^and_result12[43]^and_result12[44]^and_result12[45]^and_result12[46]^and_result12[47]^and_result12[48]^and_result12[49]^and_result12[50]^and_result12[51]^and_result12[52]^and_result12[53]^and_result12[54]^and_result12[55]^and_result12[56]^and_result12[57]^and_result12[58]^and_result12[59]^and_result12[60]^and_result12[61]^and_result12[62]^and_result12[63]^and_result12[64]^and_result12[65]^and_result12[66]^and_result12[67]^and_result12[68]^and_result12[69]^and_result12[70]^and_result12[71]^and_result12[72]^and_result12[73]^and_result12[74]^and_result12[75]^and_result12[76]^and_result12[77]^and_result12[78]^and_result12[79]^and_result12[80]^and_result12[81]^and_result12[82]^and_result12[83]^and_result12[84]^and_result12[85]^and_result12[86]^and_result12[87]^and_result12[88]^and_result12[89]^and_result12[90]^and_result12[91]^and_result12[92]^and_result12[93]^and_result12[94]^and_result12[95]^and_result12[96]^and_result12[97]^and_result12[98]^and_result12[99]^and_result12[100]^and_result12[101]^and_result12[102]^and_result12[103]^and_result12[104]^and_result12[105]^and_result12[106]^and_result12[107]^and_result12[108]^and_result12[109]^and_result12[110]^and_result12[111]^and_result12[112]^and_result12[113]^and_result12[114]^and_result12[115]^and_result12[116]^and_result12[117]^and_result12[118]^and_result12[119]^and_result12[120]^and_result12[121]^and_result12[122]^and_result12[123]^and_result12[124]^and_result12[125]^and_result12[126]^and_result12[127]^and_result12[128]^and_result12[129]^and_result12[130]^and_result12[131]^and_result12[132]^and_result12[133]^and_result12[134]^and_result12[135]^and_result12[136]^and_result12[137]^and_result12[138]^and_result12[139]^and_result12[140]^and_result12[141]^and_result12[142]^and_result12[143]^and_result12[144]^and_result12[145]^and_result12[146]^and_result12[147]^and_result12[148]^and_result12[149]^and_result12[150]^and_result12[151]^and_result12[152]^and_result12[153]^and_result12[154]^and_result12[155]^and_result12[156]^and_result12[157]^and_result12[158]^and_result12[159]^and_result12[160]^and_result12[161]^and_result12[162]^and_result12[163]^and_result12[164]^and_result12[165]^and_result12[166]^and_result12[167]^and_result12[168]^and_result12[169]^and_result12[170]^and_result12[171]^and_result12[172]^and_result12[173]^and_result12[174]^and_result12[175]^and_result12[176]^and_result12[177]^and_result12[178]^and_result12[179]^and_result12[180]^and_result12[181]^and_result12[182]^and_result12[183]^and_result12[184]^and_result12[185]^and_result12[186]^and_result12[187]^and_result12[188]^and_result12[189]^and_result12[190]^and_result12[191]^and_result12[192]^and_result12[193]^and_result12[194]^and_result12[195]^and_result12[196]^and_result12[197]^and_result12[198]^and_result12[199]^and_result12[200]^and_result12[201]^and_result12[202]^and_result12[203]^and_result12[204]^and_result12[205]^and_result12[206]^and_result12[207]^and_result12[208]^and_result12[209]^and_result12[210]^and_result12[211]^and_result12[212]^and_result12[213]^and_result12[214]^and_result12[215]^and_result12[216]^and_result12[217]^and_result12[218]^and_result12[219]^and_result12[220]^and_result12[221]^and_result12[222]^and_result12[223]^and_result12[224]^and_result12[225]^and_result12[226]^and_result12[227]^and_result12[228]^and_result12[229]^and_result12[230]^and_result12[231]^and_result12[232]^and_result12[233]^and_result12[234]^and_result12[235]^and_result12[236]^and_result12[237]^and_result12[238]^and_result12[239]^and_result12[240]^and_result12[241]^and_result12[242]^and_result12[243]^and_result12[244]^and_result12[245]^and_result12[246]^and_result12[247]^and_result12[248]^and_result12[249]^and_result12[250]^and_result12[251]^and_result12[252]^and_result12[253]^and_result12[254];
assign key[13]=and_result13[0]^and_result13[1]^and_result13[2]^and_result13[3]^and_result13[4]^and_result13[5]^and_result13[6]^and_result13[7]^and_result13[8]^and_result13[9]^and_result13[10]^and_result13[11]^and_result13[12]^and_result13[13]^and_result13[14]^and_result13[15]^and_result13[16]^and_result13[17]^and_result13[18]^and_result13[19]^and_result13[20]^and_result13[21]^and_result13[22]^and_result13[23]^and_result13[24]^and_result13[25]^and_result13[26]^and_result13[27]^and_result13[28]^and_result13[29]^and_result13[30]^and_result13[31]^and_result13[32]^and_result13[33]^and_result13[34]^and_result13[35]^and_result13[36]^and_result13[37]^and_result13[38]^and_result13[39]^and_result13[40]^and_result13[41]^and_result13[42]^and_result13[43]^and_result13[44]^and_result13[45]^and_result13[46]^and_result13[47]^and_result13[48]^and_result13[49]^and_result13[50]^and_result13[51]^and_result13[52]^and_result13[53]^and_result13[54]^and_result13[55]^and_result13[56]^and_result13[57]^and_result13[58]^and_result13[59]^and_result13[60]^and_result13[61]^and_result13[62]^and_result13[63]^and_result13[64]^and_result13[65]^and_result13[66]^and_result13[67]^and_result13[68]^and_result13[69]^and_result13[70]^and_result13[71]^and_result13[72]^and_result13[73]^and_result13[74]^and_result13[75]^and_result13[76]^and_result13[77]^and_result13[78]^and_result13[79]^and_result13[80]^and_result13[81]^and_result13[82]^and_result13[83]^and_result13[84]^and_result13[85]^and_result13[86]^and_result13[87]^and_result13[88]^and_result13[89]^and_result13[90]^and_result13[91]^and_result13[92]^and_result13[93]^and_result13[94]^and_result13[95]^and_result13[96]^and_result13[97]^and_result13[98]^and_result13[99]^and_result13[100]^and_result13[101]^and_result13[102]^and_result13[103]^and_result13[104]^and_result13[105]^and_result13[106]^and_result13[107]^and_result13[108]^and_result13[109]^and_result13[110]^and_result13[111]^and_result13[112]^and_result13[113]^and_result13[114]^and_result13[115]^and_result13[116]^and_result13[117]^and_result13[118]^and_result13[119]^and_result13[120]^and_result13[121]^and_result13[122]^and_result13[123]^and_result13[124]^and_result13[125]^and_result13[126]^and_result13[127]^and_result13[128]^and_result13[129]^and_result13[130]^and_result13[131]^and_result13[132]^and_result13[133]^and_result13[134]^and_result13[135]^and_result13[136]^and_result13[137]^and_result13[138]^and_result13[139]^and_result13[140]^and_result13[141]^and_result13[142]^and_result13[143]^and_result13[144]^and_result13[145]^and_result13[146]^and_result13[147]^and_result13[148]^and_result13[149]^and_result13[150]^and_result13[151]^and_result13[152]^and_result13[153]^and_result13[154]^and_result13[155]^and_result13[156]^and_result13[157]^and_result13[158]^and_result13[159]^and_result13[160]^and_result13[161]^and_result13[162]^and_result13[163]^and_result13[164]^and_result13[165]^and_result13[166]^and_result13[167]^and_result13[168]^and_result13[169]^and_result13[170]^and_result13[171]^and_result13[172]^and_result13[173]^and_result13[174]^and_result13[175]^and_result13[176]^and_result13[177]^and_result13[178]^and_result13[179]^and_result13[180]^and_result13[181]^and_result13[182]^and_result13[183]^and_result13[184]^and_result13[185]^and_result13[186]^and_result13[187]^and_result13[188]^and_result13[189]^and_result13[190]^and_result13[191]^and_result13[192]^and_result13[193]^and_result13[194]^and_result13[195]^and_result13[196]^and_result13[197]^and_result13[198]^and_result13[199]^and_result13[200]^and_result13[201]^and_result13[202]^and_result13[203]^and_result13[204]^and_result13[205]^and_result13[206]^and_result13[207]^and_result13[208]^and_result13[209]^and_result13[210]^and_result13[211]^and_result13[212]^and_result13[213]^and_result13[214]^and_result13[215]^and_result13[216]^and_result13[217]^and_result13[218]^and_result13[219]^and_result13[220]^and_result13[221]^and_result13[222]^and_result13[223]^and_result13[224]^and_result13[225]^and_result13[226]^and_result13[227]^and_result13[228]^and_result13[229]^and_result13[230]^and_result13[231]^and_result13[232]^and_result13[233]^and_result13[234]^and_result13[235]^and_result13[236]^and_result13[237]^and_result13[238]^and_result13[239]^and_result13[240]^and_result13[241]^and_result13[242]^and_result13[243]^and_result13[244]^and_result13[245]^and_result13[246]^and_result13[247]^and_result13[248]^and_result13[249]^and_result13[250]^and_result13[251]^and_result13[252]^and_result13[253]^and_result13[254];
assign key[14]=and_result14[0]^and_result14[1]^and_result14[2]^and_result14[3]^and_result14[4]^and_result14[5]^and_result14[6]^and_result14[7]^and_result14[8]^and_result14[9]^and_result14[10]^and_result14[11]^and_result14[12]^and_result14[13]^and_result14[14]^and_result14[15]^and_result14[16]^and_result14[17]^and_result14[18]^and_result14[19]^and_result14[20]^and_result14[21]^and_result14[22]^and_result14[23]^and_result14[24]^and_result14[25]^and_result14[26]^and_result14[27]^and_result14[28]^and_result14[29]^and_result14[30]^and_result14[31]^and_result14[32]^and_result14[33]^and_result14[34]^and_result14[35]^and_result14[36]^and_result14[37]^and_result14[38]^and_result14[39]^and_result14[40]^and_result14[41]^and_result14[42]^and_result14[43]^and_result14[44]^and_result14[45]^and_result14[46]^and_result14[47]^and_result14[48]^and_result14[49]^and_result14[50]^and_result14[51]^and_result14[52]^and_result14[53]^and_result14[54]^and_result14[55]^and_result14[56]^and_result14[57]^and_result14[58]^and_result14[59]^and_result14[60]^and_result14[61]^and_result14[62]^and_result14[63]^and_result14[64]^and_result14[65]^and_result14[66]^and_result14[67]^and_result14[68]^and_result14[69]^and_result14[70]^and_result14[71]^and_result14[72]^and_result14[73]^and_result14[74]^and_result14[75]^and_result14[76]^and_result14[77]^and_result14[78]^and_result14[79]^and_result14[80]^and_result14[81]^and_result14[82]^and_result14[83]^and_result14[84]^and_result14[85]^and_result14[86]^and_result14[87]^and_result14[88]^and_result14[89]^and_result14[90]^and_result14[91]^and_result14[92]^and_result14[93]^and_result14[94]^and_result14[95]^and_result14[96]^and_result14[97]^and_result14[98]^and_result14[99]^and_result14[100]^and_result14[101]^and_result14[102]^and_result14[103]^and_result14[104]^and_result14[105]^and_result14[106]^and_result14[107]^and_result14[108]^and_result14[109]^and_result14[110]^and_result14[111]^and_result14[112]^and_result14[113]^and_result14[114]^and_result14[115]^and_result14[116]^and_result14[117]^and_result14[118]^and_result14[119]^and_result14[120]^and_result14[121]^and_result14[122]^and_result14[123]^and_result14[124]^and_result14[125]^and_result14[126]^and_result14[127]^and_result14[128]^and_result14[129]^and_result14[130]^and_result14[131]^and_result14[132]^and_result14[133]^and_result14[134]^and_result14[135]^and_result14[136]^and_result14[137]^and_result14[138]^and_result14[139]^and_result14[140]^and_result14[141]^and_result14[142]^and_result14[143]^and_result14[144]^and_result14[145]^and_result14[146]^and_result14[147]^and_result14[148]^and_result14[149]^and_result14[150]^and_result14[151]^and_result14[152]^and_result14[153]^and_result14[154]^and_result14[155]^and_result14[156]^and_result14[157]^and_result14[158]^and_result14[159]^and_result14[160]^and_result14[161]^and_result14[162]^and_result14[163]^and_result14[164]^and_result14[165]^and_result14[166]^and_result14[167]^and_result14[168]^and_result14[169]^and_result14[170]^and_result14[171]^and_result14[172]^and_result14[173]^and_result14[174]^and_result14[175]^and_result14[176]^and_result14[177]^and_result14[178]^and_result14[179]^and_result14[180]^and_result14[181]^and_result14[182]^and_result14[183]^and_result14[184]^and_result14[185]^and_result14[186]^and_result14[187]^and_result14[188]^and_result14[189]^and_result14[190]^and_result14[191]^and_result14[192]^and_result14[193]^and_result14[194]^and_result14[195]^and_result14[196]^and_result14[197]^and_result14[198]^and_result14[199]^and_result14[200]^and_result14[201]^and_result14[202]^and_result14[203]^and_result14[204]^and_result14[205]^and_result14[206]^and_result14[207]^and_result14[208]^and_result14[209]^and_result14[210]^and_result14[211]^and_result14[212]^and_result14[213]^and_result14[214]^and_result14[215]^and_result14[216]^and_result14[217]^and_result14[218]^and_result14[219]^and_result14[220]^and_result14[221]^and_result14[222]^and_result14[223]^and_result14[224]^and_result14[225]^and_result14[226]^and_result14[227]^and_result14[228]^and_result14[229]^and_result14[230]^and_result14[231]^and_result14[232]^and_result14[233]^and_result14[234]^and_result14[235]^and_result14[236]^and_result14[237]^and_result14[238]^and_result14[239]^and_result14[240]^and_result14[241]^and_result14[242]^and_result14[243]^and_result14[244]^and_result14[245]^and_result14[246]^and_result14[247]^and_result14[248]^and_result14[249]^and_result14[250]^and_result14[251]^and_result14[252]^and_result14[253]^and_result14[254];
assign key[15]=and_result15[0]^and_result15[1]^and_result15[2]^and_result15[3]^and_result15[4]^and_result15[5]^and_result15[6]^and_result15[7]^and_result15[8]^and_result15[9]^and_result15[10]^and_result15[11]^and_result15[12]^and_result15[13]^and_result15[14]^and_result15[15]^and_result15[16]^and_result15[17]^and_result15[18]^and_result15[19]^and_result15[20]^and_result15[21]^and_result15[22]^and_result15[23]^and_result15[24]^and_result15[25]^and_result15[26]^and_result15[27]^and_result15[28]^and_result15[29]^and_result15[30]^and_result15[31]^and_result15[32]^and_result15[33]^and_result15[34]^and_result15[35]^and_result15[36]^and_result15[37]^and_result15[38]^and_result15[39]^and_result15[40]^and_result15[41]^and_result15[42]^and_result15[43]^and_result15[44]^and_result15[45]^and_result15[46]^and_result15[47]^and_result15[48]^and_result15[49]^and_result15[50]^and_result15[51]^and_result15[52]^and_result15[53]^and_result15[54]^and_result15[55]^and_result15[56]^and_result15[57]^and_result15[58]^and_result15[59]^and_result15[60]^and_result15[61]^and_result15[62]^and_result15[63]^and_result15[64]^and_result15[65]^and_result15[66]^and_result15[67]^and_result15[68]^and_result15[69]^and_result15[70]^and_result15[71]^and_result15[72]^and_result15[73]^and_result15[74]^and_result15[75]^and_result15[76]^and_result15[77]^and_result15[78]^and_result15[79]^and_result15[80]^and_result15[81]^and_result15[82]^and_result15[83]^and_result15[84]^and_result15[85]^and_result15[86]^and_result15[87]^and_result15[88]^and_result15[89]^and_result15[90]^and_result15[91]^and_result15[92]^and_result15[93]^and_result15[94]^and_result15[95]^and_result15[96]^and_result15[97]^and_result15[98]^and_result15[99]^and_result15[100]^and_result15[101]^and_result15[102]^and_result15[103]^and_result15[104]^and_result15[105]^and_result15[106]^and_result15[107]^and_result15[108]^and_result15[109]^and_result15[110]^and_result15[111]^and_result15[112]^and_result15[113]^and_result15[114]^and_result15[115]^and_result15[116]^and_result15[117]^and_result15[118]^and_result15[119]^and_result15[120]^and_result15[121]^and_result15[122]^and_result15[123]^and_result15[124]^and_result15[125]^and_result15[126]^and_result15[127]^and_result15[128]^and_result15[129]^and_result15[130]^and_result15[131]^and_result15[132]^and_result15[133]^and_result15[134]^and_result15[135]^and_result15[136]^and_result15[137]^and_result15[138]^and_result15[139]^and_result15[140]^and_result15[141]^and_result15[142]^and_result15[143]^and_result15[144]^and_result15[145]^and_result15[146]^and_result15[147]^and_result15[148]^and_result15[149]^and_result15[150]^and_result15[151]^and_result15[152]^and_result15[153]^and_result15[154]^and_result15[155]^and_result15[156]^and_result15[157]^and_result15[158]^and_result15[159]^and_result15[160]^and_result15[161]^and_result15[162]^and_result15[163]^and_result15[164]^and_result15[165]^and_result15[166]^and_result15[167]^and_result15[168]^and_result15[169]^and_result15[170]^and_result15[171]^and_result15[172]^and_result15[173]^and_result15[174]^and_result15[175]^and_result15[176]^and_result15[177]^and_result15[178]^and_result15[179]^and_result15[180]^and_result15[181]^and_result15[182]^and_result15[183]^and_result15[184]^and_result15[185]^and_result15[186]^and_result15[187]^and_result15[188]^and_result15[189]^and_result15[190]^and_result15[191]^and_result15[192]^and_result15[193]^and_result15[194]^and_result15[195]^and_result15[196]^and_result15[197]^and_result15[198]^and_result15[199]^and_result15[200]^and_result15[201]^and_result15[202]^and_result15[203]^and_result15[204]^and_result15[205]^and_result15[206]^and_result15[207]^and_result15[208]^and_result15[209]^and_result15[210]^and_result15[211]^and_result15[212]^and_result15[213]^and_result15[214]^and_result15[215]^and_result15[216]^and_result15[217]^and_result15[218]^and_result15[219]^and_result15[220]^and_result15[221]^and_result15[222]^and_result15[223]^and_result15[224]^and_result15[225]^and_result15[226]^and_result15[227]^and_result15[228]^and_result15[229]^and_result15[230]^and_result15[231]^and_result15[232]^and_result15[233]^and_result15[234]^and_result15[235]^and_result15[236]^and_result15[237]^and_result15[238]^and_result15[239]^and_result15[240]^and_result15[241]^and_result15[242]^and_result15[243]^and_result15[244]^and_result15[245]^and_result15[246]^and_result15[247]^and_result15[248]^and_result15[249]^and_result15[250]^and_result15[251]^and_result15[252]^and_result15[253]^and_result15[254];
assign key[16]=and_result16[0]^and_result16[1]^and_result16[2]^and_result16[3]^and_result16[4]^and_result16[5]^and_result16[6]^and_result16[7]^and_result16[8]^and_result16[9]^and_result16[10]^and_result16[11]^and_result16[12]^and_result16[13]^and_result16[14]^and_result16[15]^and_result16[16]^and_result16[17]^and_result16[18]^and_result16[19]^and_result16[20]^and_result16[21]^and_result16[22]^and_result16[23]^and_result16[24]^and_result16[25]^and_result16[26]^and_result16[27]^and_result16[28]^and_result16[29]^and_result16[30]^and_result16[31]^and_result16[32]^and_result16[33]^and_result16[34]^and_result16[35]^and_result16[36]^and_result16[37]^and_result16[38]^and_result16[39]^and_result16[40]^and_result16[41]^and_result16[42]^and_result16[43]^and_result16[44]^and_result16[45]^and_result16[46]^and_result16[47]^and_result16[48]^and_result16[49]^and_result16[50]^and_result16[51]^and_result16[52]^and_result16[53]^and_result16[54]^and_result16[55]^and_result16[56]^and_result16[57]^and_result16[58]^and_result16[59]^and_result16[60]^and_result16[61]^and_result16[62]^and_result16[63]^and_result16[64]^and_result16[65]^and_result16[66]^and_result16[67]^and_result16[68]^and_result16[69]^and_result16[70]^and_result16[71]^and_result16[72]^and_result16[73]^and_result16[74]^and_result16[75]^and_result16[76]^and_result16[77]^and_result16[78]^and_result16[79]^and_result16[80]^and_result16[81]^and_result16[82]^and_result16[83]^and_result16[84]^and_result16[85]^and_result16[86]^and_result16[87]^and_result16[88]^and_result16[89]^and_result16[90]^and_result16[91]^and_result16[92]^and_result16[93]^and_result16[94]^and_result16[95]^and_result16[96]^and_result16[97]^and_result16[98]^and_result16[99]^and_result16[100]^and_result16[101]^and_result16[102]^and_result16[103]^and_result16[104]^and_result16[105]^and_result16[106]^and_result16[107]^and_result16[108]^and_result16[109]^and_result16[110]^and_result16[111]^and_result16[112]^and_result16[113]^and_result16[114]^and_result16[115]^and_result16[116]^and_result16[117]^and_result16[118]^and_result16[119]^and_result16[120]^and_result16[121]^and_result16[122]^and_result16[123]^and_result16[124]^and_result16[125]^and_result16[126]^and_result16[127]^and_result16[128]^and_result16[129]^and_result16[130]^and_result16[131]^and_result16[132]^and_result16[133]^and_result16[134]^and_result16[135]^and_result16[136]^and_result16[137]^and_result16[138]^and_result16[139]^and_result16[140]^and_result16[141]^and_result16[142]^and_result16[143]^and_result16[144]^and_result16[145]^and_result16[146]^and_result16[147]^and_result16[148]^and_result16[149]^and_result16[150]^and_result16[151]^and_result16[152]^and_result16[153]^and_result16[154]^and_result16[155]^and_result16[156]^and_result16[157]^and_result16[158]^and_result16[159]^and_result16[160]^and_result16[161]^and_result16[162]^and_result16[163]^and_result16[164]^and_result16[165]^and_result16[166]^and_result16[167]^and_result16[168]^and_result16[169]^and_result16[170]^and_result16[171]^and_result16[172]^and_result16[173]^and_result16[174]^and_result16[175]^and_result16[176]^and_result16[177]^and_result16[178]^and_result16[179]^and_result16[180]^and_result16[181]^and_result16[182]^and_result16[183]^and_result16[184]^and_result16[185]^and_result16[186]^and_result16[187]^and_result16[188]^and_result16[189]^and_result16[190]^and_result16[191]^and_result16[192]^and_result16[193]^and_result16[194]^and_result16[195]^and_result16[196]^and_result16[197]^and_result16[198]^and_result16[199]^and_result16[200]^and_result16[201]^and_result16[202]^and_result16[203]^and_result16[204]^and_result16[205]^and_result16[206]^and_result16[207]^and_result16[208]^and_result16[209]^and_result16[210]^and_result16[211]^and_result16[212]^and_result16[213]^and_result16[214]^and_result16[215]^and_result16[216]^and_result16[217]^and_result16[218]^and_result16[219]^and_result16[220]^and_result16[221]^and_result16[222]^and_result16[223]^and_result16[224]^and_result16[225]^and_result16[226]^and_result16[227]^and_result16[228]^and_result16[229]^and_result16[230]^and_result16[231]^and_result16[232]^and_result16[233]^and_result16[234]^and_result16[235]^and_result16[236]^and_result16[237]^and_result16[238]^and_result16[239]^and_result16[240]^and_result16[241]^and_result16[242]^and_result16[243]^and_result16[244]^and_result16[245]^and_result16[246]^and_result16[247]^and_result16[248]^and_result16[249]^and_result16[250]^and_result16[251]^and_result16[252]^and_result16[253]^and_result16[254];
assign key[17]=and_result17[0]^and_result17[1]^and_result17[2]^and_result17[3]^and_result17[4]^and_result17[5]^and_result17[6]^and_result17[7]^and_result17[8]^and_result17[9]^and_result17[10]^and_result17[11]^and_result17[12]^and_result17[13]^and_result17[14]^and_result17[15]^and_result17[16]^and_result17[17]^and_result17[18]^and_result17[19]^and_result17[20]^and_result17[21]^and_result17[22]^and_result17[23]^and_result17[24]^and_result17[25]^and_result17[26]^and_result17[27]^and_result17[28]^and_result17[29]^and_result17[30]^and_result17[31]^and_result17[32]^and_result17[33]^and_result17[34]^and_result17[35]^and_result17[36]^and_result17[37]^and_result17[38]^and_result17[39]^and_result17[40]^and_result17[41]^and_result17[42]^and_result17[43]^and_result17[44]^and_result17[45]^and_result17[46]^and_result17[47]^and_result17[48]^and_result17[49]^and_result17[50]^and_result17[51]^and_result17[52]^and_result17[53]^and_result17[54]^and_result17[55]^and_result17[56]^and_result17[57]^and_result17[58]^and_result17[59]^and_result17[60]^and_result17[61]^and_result17[62]^and_result17[63]^and_result17[64]^and_result17[65]^and_result17[66]^and_result17[67]^and_result17[68]^and_result17[69]^and_result17[70]^and_result17[71]^and_result17[72]^and_result17[73]^and_result17[74]^and_result17[75]^and_result17[76]^and_result17[77]^and_result17[78]^and_result17[79]^and_result17[80]^and_result17[81]^and_result17[82]^and_result17[83]^and_result17[84]^and_result17[85]^and_result17[86]^and_result17[87]^and_result17[88]^and_result17[89]^and_result17[90]^and_result17[91]^and_result17[92]^and_result17[93]^and_result17[94]^and_result17[95]^and_result17[96]^and_result17[97]^and_result17[98]^and_result17[99]^and_result17[100]^and_result17[101]^and_result17[102]^and_result17[103]^and_result17[104]^and_result17[105]^and_result17[106]^and_result17[107]^and_result17[108]^and_result17[109]^and_result17[110]^and_result17[111]^and_result17[112]^and_result17[113]^and_result17[114]^and_result17[115]^and_result17[116]^and_result17[117]^and_result17[118]^and_result17[119]^and_result17[120]^and_result17[121]^and_result17[122]^and_result17[123]^and_result17[124]^and_result17[125]^and_result17[126]^and_result17[127]^and_result17[128]^and_result17[129]^and_result17[130]^and_result17[131]^and_result17[132]^and_result17[133]^and_result17[134]^and_result17[135]^and_result17[136]^and_result17[137]^and_result17[138]^and_result17[139]^and_result17[140]^and_result17[141]^and_result17[142]^and_result17[143]^and_result17[144]^and_result17[145]^and_result17[146]^and_result17[147]^and_result17[148]^and_result17[149]^and_result17[150]^and_result17[151]^and_result17[152]^and_result17[153]^and_result17[154]^and_result17[155]^and_result17[156]^and_result17[157]^and_result17[158]^and_result17[159]^and_result17[160]^and_result17[161]^and_result17[162]^and_result17[163]^and_result17[164]^and_result17[165]^and_result17[166]^and_result17[167]^and_result17[168]^and_result17[169]^and_result17[170]^and_result17[171]^and_result17[172]^and_result17[173]^and_result17[174]^and_result17[175]^and_result17[176]^and_result17[177]^and_result17[178]^and_result17[179]^and_result17[180]^and_result17[181]^and_result17[182]^and_result17[183]^and_result17[184]^and_result17[185]^and_result17[186]^and_result17[187]^and_result17[188]^and_result17[189]^and_result17[190]^and_result17[191]^and_result17[192]^and_result17[193]^and_result17[194]^and_result17[195]^and_result17[196]^and_result17[197]^and_result17[198]^and_result17[199]^and_result17[200]^and_result17[201]^and_result17[202]^and_result17[203]^and_result17[204]^and_result17[205]^and_result17[206]^and_result17[207]^and_result17[208]^and_result17[209]^and_result17[210]^and_result17[211]^and_result17[212]^and_result17[213]^and_result17[214]^and_result17[215]^and_result17[216]^and_result17[217]^and_result17[218]^and_result17[219]^and_result17[220]^and_result17[221]^and_result17[222]^and_result17[223]^and_result17[224]^and_result17[225]^and_result17[226]^and_result17[227]^and_result17[228]^and_result17[229]^and_result17[230]^and_result17[231]^and_result17[232]^and_result17[233]^and_result17[234]^and_result17[235]^and_result17[236]^and_result17[237]^and_result17[238]^and_result17[239]^and_result17[240]^and_result17[241]^and_result17[242]^and_result17[243]^and_result17[244]^and_result17[245]^and_result17[246]^and_result17[247]^and_result17[248]^and_result17[249]^and_result17[250]^and_result17[251]^and_result17[252]^and_result17[253]^and_result17[254];
assign key[18]=and_result18[0]^and_result18[1]^and_result18[2]^and_result18[3]^and_result18[4]^and_result18[5]^and_result18[6]^and_result18[7]^and_result18[8]^and_result18[9]^and_result18[10]^and_result18[11]^and_result18[12]^and_result18[13]^and_result18[14]^and_result18[15]^and_result18[16]^and_result18[17]^and_result18[18]^and_result18[19]^and_result18[20]^and_result18[21]^and_result18[22]^and_result18[23]^and_result18[24]^and_result18[25]^and_result18[26]^and_result18[27]^and_result18[28]^and_result18[29]^and_result18[30]^and_result18[31]^and_result18[32]^and_result18[33]^and_result18[34]^and_result18[35]^and_result18[36]^and_result18[37]^and_result18[38]^and_result18[39]^and_result18[40]^and_result18[41]^and_result18[42]^and_result18[43]^and_result18[44]^and_result18[45]^and_result18[46]^and_result18[47]^and_result18[48]^and_result18[49]^and_result18[50]^and_result18[51]^and_result18[52]^and_result18[53]^and_result18[54]^and_result18[55]^and_result18[56]^and_result18[57]^and_result18[58]^and_result18[59]^and_result18[60]^and_result18[61]^and_result18[62]^and_result18[63]^and_result18[64]^and_result18[65]^and_result18[66]^and_result18[67]^and_result18[68]^and_result18[69]^and_result18[70]^and_result18[71]^and_result18[72]^and_result18[73]^and_result18[74]^and_result18[75]^and_result18[76]^and_result18[77]^and_result18[78]^and_result18[79]^and_result18[80]^and_result18[81]^and_result18[82]^and_result18[83]^and_result18[84]^and_result18[85]^and_result18[86]^and_result18[87]^and_result18[88]^and_result18[89]^and_result18[90]^and_result18[91]^and_result18[92]^and_result18[93]^and_result18[94]^and_result18[95]^and_result18[96]^and_result18[97]^and_result18[98]^and_result18[99]^and_result18[100]^and_result18[101]^and_result18[102]^and_result18[103]^and_result18[104]^and_result18[105]^and_result18[106]^and_result18[107]^and_result18[108]^and_result18[109]^and_result18[110]^and_result18[111]^and_result18[112]^and_result18[113]^and_result18[114]^and_result18[115]^and_result18[116]^and_result18[117]^and_result18[118]^and_result18[119]^and_result18[120]^and_result18[121]^and_result18[122]^and_result18[123]^and_result18[124]^and_result18[125]^and_result18[126]^and_result18[127]^and_result18[128]^and_result18[129]^and_result18[130]^and_result18[131]^and_result18[132]^and_result18[133]^and_result18[134]^and_result18[135]^and_result18[136]^and_result18[137]^and_result18[138]^and_result18[139]^and_result18[140]^and_result18[141]^and_result18[142]^and_result18[143]^and_result18[144]^and_result18[145]^and_result18[146]^and_result18[147]^and_result18[148]^and_result18[149]^and_result18[150]^and_result18[151]^and_result18[152]^and_result18[153]^and_result18[154]^and_result18[155]^and_result18[156]^and_result18[157]^and_result18[158]^and_result18[159]^and_result18[160]^and_result18[161]^and_result18[162]^and_result18[163]^and_result18[164]^and_result18[165]^and_result18[166]^and_result18[167]^and_result18[168]^and_result18[169]^and_result18[170]^and_result18[171]^and_result18[172]^and_result18[173]^and_result18[174]^and_result18[175]^and_result18[176]^and_result18[177]^and_result18[178]^and_result18[179]^and_result18[180]^and_result18[181]^and_result18[182]^and_result18[183]^and_result18[184]^and_result18[185]^and_result18[186]^and_result18[187]^and_result18[188]^and_result18[189]^and_result18[190]^and_result18[191]^and_result18[192]^and_result18[193]^and_result18[194]^and_result18[195]^and_result18[196]^and_result18[197]^and_result18[198]^and_result18[199]^and_result18[200]^and_result18[201]^and_result18[202]^and_result18[203]^and_result18[204]^and_result18[205]^and_result18[206]^and_result18[207]^and_result18[208]^and_result18[209]^and_result18[210]^and_result18[211]^and_result18[212]^and_result18[213]^and_result18[214]^and_result18[215]^and_result18[216]^and_result18[217]^and_result18[218]^and_result18[219]^and_result18[220]^and_result18[221]^and_result18[222]^and_result18[223]^and_result18[224]^and_result18[225]^and_result18[226]^and_result18[227]^and_result18[228]^and_result18[229]^and_result18[230]^and_result18[231]^and_result18[232]^and_result18[233]^and_result18[234]^and_result18[235]^and_result18[236]^and_result18[237]^and_result18[238]^and_result18[239]^and_result18[240]^and_result18[241]^and_result18[242]^and_result18[243]^and_result18[244]^and_result18[245]^and_result18[246]^and_result18[247]^and_result18[248]^and_result18[249]^and_result18[250]^and_result18[251]^and_result18[252]^and_result18[253]^and_result18[254];
assign key[19]=and_result19[0]^and_result19[1]^and_result19[2]^and_result19[3]^and_result19[4]^and_result19[5]^and_result19[6]^and_result19[7]^and_result19[8]^and_result19[9]^and_result19[10]^and_result19[11]^and_result19[12]^and_result19[13]^and_result19[14]^and_result19[15]^and_result19[16]^and_result19[17]^and_result19[18]^and_result19[19]^and_result19[20]^and_result19[21]^and_result19[22]^and_result19[23]^and_result19[24]^and_result19[25]^and_result19[26]^and_result19[27]^and_result19[28]^and_result19[29]^and_result19[30]^and_result19[31]^and_result19[32]^and_result19[33]^and_result19[34]^and_result19[35]^and_result19[36]^and_result19[37]^and_result19[38]^and_result19[39]^and_result19[40]^and_result19[41]^and_result19[42]^and_result19[43]^and_result19[44]^and_result19[45]^and_result19[46]^and_result19[47]^and_result19[48]^and_result19[49]^and_result19[50]^and_result19[51]^and_result19[52]^and_result19[53]^and_result19[54]^and_result19[55]^and_result19[56]^and_result19[57]^and_result19[58]^and_result19[59]^and_result19[60]^and_result19[61]^and_result19[62]^and_result19[63]^and_result19[64]^and_result19[65]^and_result19[66]^and_result19[67]^and_result19[68]^and_result19[69]^and_result19[70]^and_result19[71]^and_result19[72]^and_result19[73]^and_result19[74]^and_result19[75]^and_result19[76]^and_result19[77]^and_result19[78]^and_result19[79]^and_result19[80]^and_result19[81]^and_result19[82]^and_result19[83]^and_result19[84]^and_result19[85]^and_result19[86]^and_result19[87]^and_result19[88]^and_result19[89]^and_result19[90]^and_result19[91]^and_result19[92]^and_result19[93]^and_result19[94]^and_result19[95]^and_result19[96]^and_result19[97]^and_result19[98]^and_result19[99]^and_result19[100]^and_result19[101]^and_result19[102]^and_result19[103]^and_result19[104]^and_result19[105]^and_result19[106]^and_result19[107]^and_result19[108]^and_result19[109]^and_result19[110]^and_result19[111]^and_result19[112]^and_result19[113]^and_result19[114]^and_result19[115]^and_result19[116]^and_result19[117]^and_result19[118]^and_result19[119]^and_result19[120]^and_result19[121]^and_result19[122]^and_result19[123]^and_result19[124]^and_result19[125]^and_result19[126]^and_result19[127]^and_result19[128]^and_result19[129]^and_result19[130]^and_result19[131]^and_result19[132]^and_result19[133]^and_result19[134]^and_result19[135]^and_result19[136]^and_result19[137]^and_result19[138]^and_result19[139]^and_result19[140]^and_result19[141]^and_result19[142]^and_result19[143]^and_result19[144]^and_result19[145]^and_result19[146]^and_result19[147]^and_result19[148]^and_result19[149]^and_result19[150]^and_result19[151]^and_result19[152]^and_result19[153]^and_result19[154]^and_result19[155]^and_result19[156]^and_result19[157]^and_result19[158]^and_result19[159]^and_result19[160]^and_result19[161]^and_result19[162]^and_result19[163]^and_result19[164]^and_result19[165]^and_result19[166]^and_result19[167]^and_result19[168]^and_result19[169]^and_result19[170]^and_result19[171]^and_result19[172]^and_result19[173]^and_result19[174]^and_result19[175]^and_result19[176]^and_result19[177]^and_result19[178]^and_result19[179]^and_result19[180]^and_result19[181]^and_result19[182]^and_result19[183]^and_result19[184]^and_result19[185]^and_result19[186]^and_result19[187]^and_result19[188]^and_result19[189]^and_result19[190]^and_result19[191]^and_result19[192]^and_result19[193]^and_result19[194]^and_result19[195]^and_result19[196]^and_result19[197]^and_result19[198]^and_result19[199]^and_result19[200]^and_result19[201]^and_result19[202]^and_result19[203]^and_result19[204]^and_result19[205]^and_result19[206]^and_result19[207]^and_result19[208]^and_result19[209]^and_result19[210]^and_result19[211]^and_result19[212]^and_result19[213]^and_result19[214]^and_result19[215]^and_result19[216]^and_result19[217]^and_result19[218]^and_result19[219]^and_result19[220]^and_result19[221]^and_result19[222]^and_result19[223]^and_result19[224]^and_result19[225]^and_result19[226]^and_result19[227]^and_result19[228]^and_result19[229]^and_result19[230]^and_result19[231]^and_result19[232]^and_result19[233]^and_result19[234]^and_result19[235]^and_result19[236]^and_result19[237]^and_result19[238]^and_result19[239]^and_result19[240]^and_result19[241]^and_result19[242]^and_result19[243]^and_result19[244]^and_result19[245]^and_result19[246]^and_result19[247]^and_result19[248]^and_result19[249]^and_result19[250]^and_result19[251]^and_result19[252]^and_result19[253]^and_result19[254];
assign key[20]=and_result20[0]^and_result20[1]^and_result20[2]^and_result20[3]^and_result20[4]^and_result20[5]^and_result20[6]^and_result20[7]^and_result20[8]^and_result20[9]^and_result20[10]^and_result20[11]^and_result20[12]^and_result20[13]^and_result20[14]^and_result20[15]^and_result20[16]^and_result20[17]^and_result20[18]^and_result20[19]^and_result20[20]^and_result20[21]^and_result20[22]^and_result20[23]^and_result20[24]^and_result20[25]^and_result20[26]^and_result20[27]^and_result20[28]^and_result20[29]^and_result20[30]^and_result20[31]^and_result20[32]^and_result20[33]^and_result20[34]^and_result20[35]^and_result20[36]^and_result20[37]^and_result20[38]^and_result20[39]^and_result20[40]^and_result20[41]^and_result20[42]^and_result20[43]^and_result20[44]^and_result20[45]^and_result20[46]^and_result20[47]^and_result20[48]^and_result20[49]^and_result20[50]^and_result20[51]^and_result20[52]^and_result20[53]^and_result20[54]^and_result20[55]^and_result20[56]^and_result20[57]^and_result20[58]^and_result20[59]^and_result20[60]^and_result20[61]^and_result20[62]^and_result20[63]^and_result20[64]^and_result20[65]^and_result20[66]^and_result20[67]^and_result20[68]^and_result20[69]^and_result20[70]^and_result20[71]^and_result20[72]^and_result20[73]^and_result20[74]^and_result20[75]^and_result20[76]^and_result20[77]^and_result20[78]^and_result20[79]^and_result20[80]^and_result20[81]^and_result20[82]^and_result20[83]^and_result20[84]^and_result20[85]^and_result20[86]^and_result20[87]^and_result20[88]^and_result20[89]^and_result20[90]^and_result20[91]^and_result20[92]^and_result20[93]^and_result20[94]^and_result20[95]^and_result20[96]^and_result20[97]^and_result20[98]^and_result20[99]^and_result20[100]^and_result20[101]^and_result20[102]^and_result20[103]^and_result20[104]^and_result20[105]^and_result20[106]^and_result20[107]^and_result20[108]^and_result20[109]^and_result20[110]^and_result20[111]^and_result20[112]^and_result20[113]^and_result20[114]^and_result20[115]^and_result20[116]^and_result20[117]^and_result20[118]^and_result20[119]^and_result20[120]^and_result20[121]^and_result20[122]^and_result20[123]^and_result20[124]^and_result20[125]^and_result20[126]^and_result20[127]^and_result20[128]^and_result20[129]^and_result20[130]^and_result20[131]^and_result20[132]^and_result20[133]^and_result20[134]^and_result20[135]^and_result20[136]^and_result20[137]^and_result20[138]^and_result20[139]^and_result20[140]^and_result20[141]^and_result20[142]^and_result20[143]^and_result20[144]^and_result20[145]^and_result20[146]^and_result20[147]^and_result20[148]^and_result20[149]^and_result20[150]^and_result20[151]^and_result20[152]^and_result20[153]^and_result20[154]^and_result20[155]^and_result20[156]^and_result20[157]^and_result20[158]^and_result20[159]^and_result20[160]^and_result20[161]^and_result20[162]^and_result20[163]^and_result20[164]^and_result20[165]^and_result20[166]^and_result20[167]^and_result20[168]^and_result20[169]^and_result20[170]^and_result20[171]^and_result20[172]^and_result20[173]^and_result20[174]^and_result20[175]^and_result20[176]^and_result20[177]^and_result20[178]^and_result20[179]^and_result20[180]^and_result20[181]^and_result20[182]^and_result20[183]^and_result20[184]^and_result20[185]^and_result20[186]^and_result20[187]^and_result20[188]^and_result20[189]^and_result20[190]^and_result20[191]^and_result20[192]^and_result20[193]^and_result20[194]^and_result20[195]^and_result20[196]^and_result20[197]^and_result20[198]^and_result20[199]^and_result20[200]^and_result20[201]^and_result20[202]^and_result20[203]^and_result20[204]^and_result20[205]^and_result20[206]^and_result20[207]^and_result20[208]^and_result20[209]^and_result20[210]^and_result20[211]^and_result20[212]^and_result20[213]^and_result20[214]^and_result20[215]^and_result20[216]^and_result20[217]^and_result20[218]^and_result20[219]^and_result20[220]^and_result20[221]^and_result20[222]^and_result20[223]^and_result20[224]^and_result20[225]^and_result20[226]^and_result20[227]^and_result20[228]^and_result20[229]^and_result20[230]^and_result20[231]^and_result20[232]^and_result20[233]^and_result20[234]^and_result20[235]^and_result20[236]^and_result20[237]^and_result20[238]^and_result20[239]^and_result20[240]^and_result20[241]^and_result20[242]^and_result20[243]^and_result20[244]^and_result20[245]^and_result20[246]^and_result20[247]^and_result20[248]^and_result20[249]^and_result20[250]^and_result20[251]^and_result20[252]^and_result20[253]^and_result20[254];
assign key[21]=and_result21[0]^and_result21[1]^and_result21[2]^and_result21[3]^and_result21[4]^and_result21[5]^and_result21[6]^and_result21[7]^and_result21[8]^and_result21[9]^and_result21[10]^and_result21[11]^and_result21[12]^and_result21[13]^and_result21[14]^and_result21[15]^and_result21[16]^and_result21[17]^and_result21[18]^and_result21[19]^and_result21[20]^and_result21[21]^and_result21[22]^and_result21[23]^and_result21[24]^and_result21[25]^and_result21[26]^and_result21[27]^and_result21[28]^and_result21[29]^and_result21[30]^and_result21[31]^and_result21[32]^and_result21[33]^and_result21[34]^and_result21[35]^and_result21[36]^and_result21[37]^and_result21[38]^and_result21[39]^and_result21[40]^and_result21[41]^and_result21[42]^and_result21[43]^and_result21[44]^and_result21[45]^and_result21[46]^and_result21[47]^and_result21[48]^and_result21[49]^and_result21[50]^and_result21[51]^and_result21[52]^and_result21[53]^and_result21[54]^and_result21[55]^and_result21[56]^and_result21[57]^and_result21[58]^and_result21[59]^and_result21[60]^and_result21[61]^and_result21[62]^and_result21[63]^and_result21[64]^and_result21[65]^and_result21[66]^and_result21[67]^and_result21[68]^and_result21[69]^and_result21[70]^and_result21[71]^and_result21[72]^and_result21[73]^and_result21[74]^and_result21[75]^and_result21[76]^and_result21[77]^and_result21[78]^and_result21[79]^and_result21[80]^and_result21[81]^and_result21[82]^and_result21[83]^and_result21[84]^and_result21[85]^and_result21[86]^and_result21[87]^and_result21[88]^and_result21[89]^and_result21[90]^and_result21[91]^and_result21[92]^and_result21[93]^and_result21[94]^and_result21[95]^and_result21[96]^and_result21[97]^and_result21[98]^and_result21[99]^and_result21[100]^and_result21[101]^and_result21[102]^and_result21[103]^and_result21[104]^and_result21[105]^and_result21[106]^and_result21[107]^and_result21[108]^and_result21[109]^and_result21[110]^and_result21[111]^and_result21[112]^and_result21[113]^and_result21[114]^and_result21[115]^and_result21[116]^and_result21[117]^and_result21[118]^and_result21[119]^and_result21[120]^and_result21[121]^and_result21[122]^and_result21[123]^and_result21[124]^and_result21[125]^and_result21[126]^and_result21[127]^and_result21[128]^and_result21[129]^and_result21[130]^and_result21[131]^and_result21[132]^and_result21[133]^and_result21[134]^and_result21[135]^and_result21[136]^and_result21[137]^and_result21[138]^and_result21[139]^and_result21[140]^and_result21[141]^and_result21[142]^and_result21[143]^and_result21[144]^and_result21[145]^and_result21[146]^and_result21[147]^and_result21[148]^and_result21[149]^and_result21[150]^and_result21[151]^and_result21[152]^and_result21[153]^and_result21[154]^and_result21[155]^and_result21[156]^and_result21[157]^and_result21[158]^and_result21[159]^and_result21[160]^and_result21[161]^and_result21[162]^and_result21[163]^and_result21[164]^and_result21[165]^and_result21[166]^and_result21[167]^and_result21[168]^and_result21[169]^and_result21[170]^and_result21[171]^and_result21[172]^and_result21[173]^and_result21[174]^and_result21[175]^and_result21[176]^and_result21[177]^and_result21[178]^and_result21[179]^and_result21[180]^and_result21[181]^and_result21[182]^and_result21[183]^and_result21[184]^and_result21[185]^and_result21[186]^and_result21[187]^and_result21[188]^and_result21[189]^and_result21[190]^and_result21[191]^and_result21[192]^and_result21[193]^and_result21[194]^and_result21[195]^and_result21[196]^and_result21[197]^and_result21[198]^and_result21[199]^and_result21[200]^and_result21[201]^and_result21[202]^and_result21[203]^and_result21[204]^and_result21[205]^and_result21[206]^and_result21[207]^and_result21[208]^and_result21[209]^and_result21[210]^and_result21[211]^and_result21[212]^and_result21[213]^and_result21[214]^and_result21[215]^and_result21[216]^and_result21[217]^and_result21[218]^and_result21[219]^and_result21[220]^and_result21[221]^and_result21[222]^and_result21[223]^and_result21[224]^and_result21[225]^and_result21[226]^and_result21[227]^and_result21[228]^and_result21[229]^and_result21[230]^and_result21[231]^and_result21[232]^and_result21[233]^and_result21[234]^and_result21[235]^and_result21[236]^and_result21[237]^and_result21[238]^and_result21[239]^and_result21[240]^and_result21[241]^and_result21[242]^and_result21[243]^and_result21[244]^and_result21[245]^and_result21[246]^and_result21[247]^and_result21[248]^and_result21[249]^and_result21[250]^and_result21[251]^and_result21[252]^and_result21[253]^and_result21[254];
assign key[22]=and_result22[0]^and_result22[1]^and_result22[2]^and_result22[3]^and_result22[4]^and_result22[5]^and_result22[6]^and_result22[7]^and_result22[8]^and_result22[9]^and_result22[10]^and_result22[11]^and_result22[12]^and_result22[13]^and_result22[14]^and_result22[15]^and_result22[16]^and_result22[17]^and_result22[18]^and_result22[19]^and_result22[20]^and_result22[21]^and_result22[22]^and_result22[23]^and_result22[24]^and_result22[25]^and_result22[26]^and_result22[27]^and_result22[28]^and_result22[29]^and_result22[30]^and_result22[31]^and_result22[32]^and_result22[33]^and_result22[34]^and_result22[35]^and_result22[36]^and_result22[37]^and_result22[38]^and_result22[39]^and_result22[40]^and_result22[41]^and_result22[42]^and_result22[43]^and_result22[44]^and_result22[45]^and_result22[46]^and_result22[47]^and_result22[48]^and_result22[49]^and_result22[50]^and_result22[51]^and_result22[52]^and_result22[53]^and_result22[54]^and_result22[55]^and_result22[56]^and_result22[57]^and_result22[58]^and_result22[59]^and_result22[60]^and_result22[61]^and_result22[62]^and_result22[63]^and_result22[64]^and_result22[65]^and_result22[66]^and_result22[67]^and_result22[68]^and_result22[69]^and_result22[70]^and_result22[71]^and_result22[72]^and_result22[73]^and_result22[74]^and_result22[75]^and_result22[76]^and_result22[77]^and_result22[78]^and_result22[79]^and_result22[80]^and_result22[81]^and_result22[82]^and_result22[83]^and_result22[84]^and_result22[85]^and_result22[86]^and_result22[87]^and_result22[88]^and_result22[89]^and_result22[90]^and_result22[91]^and_result22[92]^and_result22[93]^and_result22[94]^and_result22[95]^and_result22[96]^and_result22[97]^and_result22[98]^and_result22[99]^and_result22[100]^and_result22[101]^and_result22[102]^and_result22[103]^and_result22[104]^and_result22[105]^and_result22[106]^and_result22[107]^and_result22[108]^and_result22[109]^and_result22[110]^and_result22[111]^and_result22[112]^and_result22[113]^and_result22[114]^and_result22[115]^and_result22[116]^and_result22[117]^and_result22[118]^and_result22[119]^and_result22[120]^and_result22[121]^and_result22[122]^and_result22[123]^and_result22[124]^and_result22[125]^and_result22[126]^and_result22[127]^and_result22[128]^and_result22[129]^and_result22[130]^and_result22[131]^and_result22[132]^and_result22[133]^and_result22[134]^and_result22[135]^and_result22[136]^and_result22[137]^and_result22[138]^and_result22[139]^and_result22[140]^and_result22[141]^and_result22[142]^and_result22[143]^and_result22[144]^and_result22[145]^and_result22[146]^and_result22[147]^and_result22[148]^and_result22[149]^and_result22[150]^and_result22[151]^and_result22[152]^and_result22[153]^and_result22[154]^and_result22[155]^and_result22[156]^and_result22[157]^and_result22[158]^and_result22[159]^and_result22[160]^and_result22[161]^and_result22[162]^and_result22[163]^and_result22[164]^and_result22[165]^and_result22[166]^and_result22[167]^and_result22[168]^and_result22[169]^and_result22[170]^and_result22[171]^and_result22[172]^and_result22[173]^and_result22[174]^and_result22[175]^and_result22[176]^and_result22[177]^and_result22[178]^and_result22[179]^and_result22[180]^and_result22[181]^and_result22[182]^and_result22[183]^and_result22[184]^and_result22[185]^and_result22[186]^and_result22[187]^and_result22[188]^and_result22[189]^and_result22[190]^and_result22[191]^and_result22[192]^and_result22[193]^and_result22[194]^and_result22[195]^and_result22[196]^and_result22[197]^and_result22[198]^and_result22[199]^and_result22[200]^and_result22[201]^and_result22[202]^and_result22[203]^and_result22[204]^and_result22[205]^and_result22[206]^and_result22[207]^and_result22[208]^and_result22[209]^and_result22[210]^and_result22[211]^and_result22[212]^and_result22[213]^and_result22[214]^and_result22[215]^and_result22[216]^and_result22[217]^and_result22[218]^and_result22[219]^and_result22[220]^and_result22[221]^and_result22[222]^and_result22[223]^and_result22[224]^and_result22[225]^and_result22[226]^and_result22[227]^and_result22[228]^and_result22[229]^and_result22[230]^and_result22[231]^and_result22[232]^and_result22[233]^and_result22[234]^and_result22[235]^and_result22[236]^and_result22[237]^and_result22[238]^and_result22[239]^and_result22[240]^and_result22[241]^and_result22[242]^and_result22[243]^and_result22[244]^and_result22[245]^and_result22[246]^and_result22[247]^and_result22[248]^and_result22[249]^and_result22[250]^and_result22[251]^and_result22[252]^and_result22[253]^and_result22[254];
assign key[23]=and_result23[0]^and_result23[1]^and_result23[2]^and_result23[3]^and_result23[4]^and_result23[5]^and_result23[6]^and_result23[7]^and_result23[8]^and_result23[9]^and_result23[10]^and_result23[11]^and_result23[12]^and_result23[13]^and_result23[14]^and_result23[15]^and_result23[16]^and_result23[17]^and_result23[18]^and_result23[19]^and_result23[20]^and_result23[21]^and_result23[22]^and_result23[23]^and_result23[24]^and_result23[25]^and_result23[26]^and_result23[27]^and_result23[28]^and_result23[29]^and_result23[30]^and_result23[31]^and_result23[32]^and_result23[33]^and_result23[34]^and_result23[35]^and_result23[36]^and_result23[37]^and_result23[38]^and_result23[39]^and_result23[40]^and_result23[41]^and_result23[42]^and_result23[43]^and_result23[44]^and_result23[45]^and_result23[46]^and_result23[47]^and_result23[48]^and_result23[49]^and_result23[50]^and_result23[51]^and_result23[52]^and_result23[53]^and_result23[54]^and_result23[55]^and_result23[56]^and_result23[57]^and_result23[58]^and_result23[59]^and_result23[60]^and_result23[61]^and_result23[62]^and_result23[63]^and_result23[64]^and_result23[65]^and_result23[66]^and_result23[67]^and_result23[68]^and_result23[69]^and_result23[70]^and_result23[71]^and_result23[72]^and_result23[73]^and_result23[74]^and_result23[75]^and_result23[76]^and_result23[77]^and_result23[78]^and_result23[79]^and_result23[80]^and_result23[81]^and_result23[82]^and_result23[83]^and_result23[84]^and_result23[85]^and_result23[86]^and_result23[87]^and_result23[88]^and_result23[89]^and_result23[90]^and_result23[91]^and_result23[92]^and_result23[93]^and_result23[94]^and_result23[95]^and_result23[96]^and_result23[97]^and_result23[98]^and_result23[99]^and_result23[100]^and_result23[101]^and_result23[102]^and_result23[103]^and_result23[104]^and_result23[105]^and_result23[106]^and_result23[107]^and_result23[108]^and_result23[109]^and_result23[110]^and_result23[111]^and_result23[112]^and_result23[113]^and_result23[114]^and_result23[115]^and_result23[116]^and_result23[117]^and_result23[118]^and_result23[119]^and_result23[120]^and_result23[121]^and_result23[122]^and_result23[123]^and_result23[124]^and_result23[125]^and_result23[126]^and_result23[127]^and_result23[128]^and_result23[129]^and_result23[130]^and_result23[131]^and_result23[132]^and_result23[133]^and_result23[134]^and_result23[135]^and_result23[136]^and_result23[137]^and_result23[138]^and_result23[139]^and_result23[140]^and_result23[141]^and_result23[142]^and_result23[143]^and_result23[144]^and_result23[145]^and_result23[146]^and_result23[147]^and_result23[148]^and_result23[149]^and_result23[150]^and_result23[151]^and_result23[152]^and_result23[153]^and_result23[154]^and_result23[155]^and_result23[156]^and_result23[157]^and_result23[158]^and_result23[159]^and_result23[160]^and_result23[161]^and_result23[162]^and_result23[163]^and_result23[164]^and_result23[165]^and_result23[166]^and_result23[167]^and_result23[168]^and_result23[169]^and_result23[170]^and_result23[171]^and_result23[172]^and_result23[173]^and_result23[174]^and_result23[175]^and_result23[176]^and_result23[177]^and_result23[178]^and_result23[179]^and_result23[180]^and_result23[181]^and_result23[182]^and_result23[183]^and_result23[184]^and_result23[185]^and_result23[186]^and_result23[187]^and_result23[188]^and_result23[189]^and_result23[190]^and_result23[191]^and_result23[192]^and_result23[193]^and_result23[194]^and_result23[195]^and_result23[196]^and_result23[197]^and_result23[198]^and_result23[199]^and_result23[200]^and_result23[201]^and_result23[202]^and_result23[203]^and_result23[204]^and_result23[205]^and_result23[206]^and_result23[207]^and_result23[208]^and_result23[209]^and_result23[210]^and_result23[211]^and_result23[212]^and_result23[213]^and_result23[214]^and_result23[215]^and_result23[216]^and_result23[217]^and_result23[218]^and_result23[219]^and_result23[220]^and_result23[221]^and_result23[222]^and_result23[223]^and_result23[224]^and_result23[225]^and_result23[226]^and_result23[227]^and_result23[228]^and_result23[229]^and_result23[230]^and_result23[231]^and_result23[232]^and_result23[233]^and_result23[234]^and_result23[235]^and_result23[236]^and_result23[237]^and_result23[238]^and_result23[239]^and_result23[240]^and_result23[241]^and_result23[242]^and_result23[243]^and_result23[244]^and_result23[245]^and_result23[246]^and_result23[247]^and_result23[248]^and_result23[249]^and_result23[250]^and_result23[251]^and_result23[252]^and_result23[253]^and_result23[254];
assign key[24]=and_result24[0]^and_result24[1]^and_result24[2]^and_result24[3]^and_result24[4]^and_result24[5]^and_result24[6]^and_result24[7]^and_result24[8]^and_result24[9]^and_result24[10]^and_result24[11]^and_result24[12]^and_result24[13]^and_result24[14]^and_result24[15]^and_result24[16]^and_result24[17]^and_result24[18]^and_result24[19]^and_result24[20]^and_result24[21]^and_result24[22]^and_result24[23]^and_result24[24]^and_result24[25]^and_result24[26]^and_result24[27]^and_result24[28]^and_result24[29]^and_result24[30]^and_result24[31]^and_result24[32]^and_result24[33]^and_result24[34]^and_result24[35]^and_result24[36]^and_result24[37]^and_result24[38]^and_result24[39]^and_result24[40]^and_result24[41]^and_result24[42]^and_result24[43]^and_result24[44]^and_result24[45]^and_result24[46]^and_result24[47]^and_result24[48]^and_result24[49]^and_result24[50]^and_result24[51]^and_result24[52]^and_result24[53]^and_result24[54]^and_result24[55]^and_result24[56]^and_result24[57]^and_result24[58]^and_result24[59]^and_result24[60]^and_result24[61]^and_result24[62]^and_result24[63]^and_result24[64]^and_result24[65]^and_result24[66]^and_result24[67]^and_result24[68]^and_result24[69]^and_result24[70]^and_result24[71]^and_result24[72]^and_result24[73]^and_result24[74]^and_result24[75]^and_result24[76]^and_result24[77]^and_result24[78]^and_result24[79]^and_result24[80]^and_result24[81]^and_result24[82]^and_result24[83]^and_result24[84]^and_result24[85]^and_result24[86]^and_result24[87]^and_result24[88]^and_result24[89]^and_result24[90]^and_result24[91]^and_result24[92]^and_result24[93]^and_result24[94]^and_result24[95]^and_result24[96]^and_result24[97]^and_result24[98]^and_result24[99]^and_result24[100]^and_result24[101]^and_result24[102]^and_result24[103]^and_result24[104]^and_result24[105]^and_result24[106]^and_result24[107]^and_result24[108]^and_result24[109]^and_result24[110]^and_result24[111]^and_result24[112]^and_result24[113]^and_result24[114]^and_result24[115]^and_result24[116]^and_result24[117]^and_result24[118]^and_result24[119]^and_result24[120]^and_result24[121]^and_result24[122]^and_result24[123]^and_result24[124]^and_result24[125]^and_result24[126]^and_result24[127]^and_result24[128]^and_result24[129]^and_result24[130]^and_result24[131]^and_result24[132]^and_result24[133]^and_result24[134]^and_result24[135]^and_result24[136]^and_result24[137]^and_result24[138]^and_result24[139]^and_result24[140]^and_result24[141]^and_result24[142]^and_result24[143]^and_result24[144]^and_result24[145]^and_result24[146]^and_result24[147]^and_result24[148]^and_result24[149]^and_result24[150]^and_result24[151]^and_result24[152]^and_result24[153]^and_result24[154]^and_result24[155]^and_result24[156]^and_result24[157]^and_result24[158]^and_result24[159]^and_result24[160]^and_result24[161]^and_result24[162]^and_result24[163]^and_result24[164]^and_result24[165]^and_result24[166]^and_result24[167]^and_result24[168]^and_result24[169]^and_result24[170]^and_result24[171]^and_result24[172]^and_result24[173]^and_result24[174]^and_result24[175]^and_result24[176]^and_result24[177]^and_result24[178]^and_result24[179]^and_result24[180]^and_result24[181]^and_result24[182]^and_result24[183]^and_result24[184]^and_result24[185]^and_result24[186]^and_result24[187]^and_result24[188]^and_result24[189]^and_result24[190]^and_result24[191]^and_result24[192]^and_result24[193]^and_result24[194]^and_result24[195]^and_result24[196]^and_result24[197]^and_result24[198]^and_result24[199]^and_result24[200]^and_result24[201]^and_result24[202]^and_result24[203]^and_result24[204]^and_result24[205]^and_result24[206]^and_result24[207]^and_result24[208]^and_result24[209]^and_result24[210]^and_result24[211]^and_result24[212]^and_result24[213]^and_result24[214]^and_result24[215]^and_result24[216]^and_result24[217]^and_result24[218]^and_result24[219]^and_result24[220]^and_result24[221]^and_result24[222]^and_result24[223]^and_result24[224]^and_result24[225]^and_result24[226]^and_result24[227]^and_result24[228]^and_result24[229]^and_result24[230]^and_result24[231]^and_result24[232]^and_result24[233]^and_result24[234]^and_result24[235]^and_result24[236]^and_result24[237]^and_result24[238]^and_result24[239]^and_result24[240]^and_result24[241]^and_result24[242]^and_result24[243]^and_result24[244]^and_result24[245]^and_result24[246]^and_result24[247]^and_result24[248]^and_result24[249]^and_result24[250]^and_result24[251]^and_result24[252]^and_result24[253]^and_result24[254];
assign key[25]=and_result25[0]^and_result25[1]^and_result25[2]^and_result25[3]^and_result25[4]^and_result25[5]^and_result25[6]^and_result25[7]^and_result25[8]^and_result25[9]^and_result25[10]^and_result25[11]^and_result25[12]^and_result25[13]^and_result25[14]^and_result25[15]^and_result25[16]^and_result25[17]^and_result25[18]^and_result25[19]^and_result25[20]^and_result25[21]^and_result25[22]^and_result25[23]^and_result25[24]^and_result25[25]^and_result25[26]^and_result25[27]^and_result25[28]^and_result25[29]^and_result25[30]^and_result25[31]^and_result25[32]^and_result25[33]^and_result25[34]^and_result25[35]^and_result25[36]^and_result25[37]^and_result25[38]^and_result25[39]^and_result25[40]^and_result25[41]^and_result25[42]^and_result25[43]^and_result25[44]^and_result25[45]^and_result25[46]^and_result25[47]^and_result25[48]^and_result25[49]^and_result25[50]^and_result25[51]^and_result25[52]^and_result25[53]^and_result25[54]^and_result25[55]^and_result25[56]^and_result25[57]^and_result25[58]^and_result25[59]^and_result25[60]^and_result25[61]^and_result25[62]^and_result25[63]^and_result25[64]^and_result25[65]^and_result25[66]^and_result25[67]^and_result25[68]^and_result25[69]^and_result25[70]^and_result25[71]^and_result25[72]^and_result25[73]^and_result25[74]^and_result25[75]^and_result25[76]^and_result25[77]^and_result25[78]^and_result25[79]^and_result25[80]^and_result25[81]^and_result25[82]^and_result25[83]^and_result25[84]^and_result25[85]^and_result25[86]^and_result25[87]^and_result25[88]^and_result25[89]^and_result25[90]^and_result25[91]^and_result25[92]^and_result25[93]^and_result25[94]^and_result25[95]^and_result25[96]^and_result25[97]^and_result25[98]^and_result25[99]^and_result25[100]^and_result25[101]^and_result25[102]^and_result25[103]^and_result25[104]^and_result25[105]^and_result25[106]^and_result25[107]^and_result25[108]^and_result25[109]^and_result25[110]^and_result25[111]^and_result25[112]^and_result25[113]^and_result25[114]^and_result25[115]^and_result25[116]^and_result25[117]^and_result25[118]^and_result25[119]^and_result25[120]^and_result25[121]^and_result25[122]^and_result25[123]^and_result25[124]^and_result25[125]^and_result25[126]^and_result25[127]^and_result25[128]^and_result25[129]^and_result25[130]^and_result25[131]^and_result25[132]^and_result25[133]^and_result25[134]^and_result25[135]^and_result25[136]^and_result25[137]^and_result25[138]^and_result25[139]^and_result25[140]^and_result25[141]^and_result25[142]^and_result25[143]^and_result25[144]^and_result25[145]^and_result25[146]^and_result25[147]^and_result25[148]^and_result25[149]^and_result25[150]^and_result25[151]^and_result25[152]^and_result25[153]^and_result25[154]^and_result25[155]^and_result25[156]^and_result25[157]^and_result25[158]^and_result25[159]^and_result25[160]^and_result25[161]^and_result25[162]^and_result25[163]^and_result25[164]^and_result25[165]^and_result25[166]^and_result25[167]^and_result25[168]^and_result25[169]^and_result25[170]^and_result25[171]^and_result25[172]^and_result25[173]^and_result25[174]^and_result25[175]^and_result25[176]^and_result25[177]^and_result25[178]^and_result25[179]^and_result25[180]^and_result25[181]^and_result25[182]^and_result25[183]^and_result25[184]^and_result25[185]^and_result25[186]^and_result25[187]^and_result25[188]^and_result25[189]^and_result25[190]^and_result25[191]^and_result25[192]^and_result25[193]^and_result25[194]^and_result25[195]^and_result25[196]^and_result25[197]^and_result25[198]^and_result25[199]^and_result25[200]^and_result25[201]^and_result25[202]^and_result25[203]^and_result25[204]^and_result25[205]^and_result25[206]^and_result25[207]^and_result25[208]^and_result25[209]^and_result25[210]^and_result25[211]^and_result25[212]^and_result25[213]^and_result25[214]^and_result25[215]^and_result25[216]^and_result25[217]^and_result25[218]^and_result25[219]^and_result25[220]^and_result25[221]^and_result25[222]^and_result25[223]^and_result25[224]^and_result25[225]^and_result25[226]^and_result25[227]^and_result25[228]^and_result25[229]^and_result25[230]^and_result25[231]^and_result25[232]^and_result25[233]^and_result25[234]^and_result25[235]^and_result25[236]^and_result25[237]^and_result25[238]^and_result25[239]^and_result25[240]^and_result25[241]^and_result25[242]^and_result25[243]^and_result25[244]^and_result25[245]^and_result25[246]^and_result25[247]^and_result25[248]^and_result25[249]^and_result25[250]^and_result25[251]^and_result25[252]^and_result25[253]^and_result25[254];
assign key[26]=and_result26[0]^and_result26[1]^and_result26[2]^and_result26[3]^and_result26[4]^and_result26[5]^and_result26[6]^and_result26[7]^and_result26[8]^and_result26[9]^and_result26[10]^and_result26[11]^and_result26[12]^and_result26[13]^and_result26[14]^and_result26[15]^and_result26[16]^and_result26[17]^and_result26[18]^and_result26[19]^and_result26[20]^and_result26[21]^and_result26[22]^and_result26[23]^and_result26[24]^and_result26[25]^and_result26[26]^and_result26[27]^and_result26[28]^and_result26[29]^and_result26[30]^and_result26[31]^and_result26[32]^and_result26[33]^and_result26[34]^and_result26[35]^and_result26[36]^and_result26[37]^and_result26[38]^and_result26[39]^and_result26[40]^and_result26[41]^and_result26[42]^and_result26[43]^and_result26[44]^and_result26[45]^and_result26[46]^and_result26[47]^and_result26[48]^and_result26[49]^and_result26[50]^and_result26[51]^and_result26[52]^and_result26[53]^and_result26[54]^and_result26[55]^and_result26[56]^and_result26[57]^and_result26[58]^and_result26[59]^and_result26[60]^and_result26[61]^and_result26[62]^and_result26[63]^and_result26[64]^and_result26[65]^and_result26[66]^and_result26[67]^and_result26[68]^and_result26[69]^and_result26[70]^and_result26[71]^and_result26[72]^and_result26[73]^and_result26[74]^and_result26[75]^and_result26[76]^and_result26[77]^and_result26[78]^and_result26[79]^and_result26[80]^and_result26[81]^and_result26[82]^and_result26[83]^and_result26[84]^and_result26[85]^and_result26[86]^and_result26[87]^and_result26[88]^and_result26[89]^and_result26[90]^and_result26[91]^and_result26[92]^and_result26[93]^and_result26[94]^and_result26[95]^and_result26[96]^and_result26[97]^and_result26[98]^and_result26[99]^and_result26[100]^and_result26[101]^and_result26[102]^and_result26[103]^and_result26[104]^and_result26[105]^and_result26[106]^and_result26[107]^and_result26[108]^and_result26[109]^and_result26[110]^and_result26[111]^and_result26[112]^and_result26[113]^and_result26[114]^and_result26[115]^and_result26[116]^and_result26[117]^and_result26[118]^and_result26[119]^and_result26[120]^and_result26[121]^and_result26[122]^and_result26[123]^and_result26[124]^and_result26[125]^and_result26[126]^and_result26[127]^and_result26[128]^and_result26[129]^and_result26[130]^and_result26[131]^and_result26[132]^and_result26[133]^and_result26[134]^and_result26[135]^and_result26[136]^and_result26[137]^and_result26[138]^and_result26[139]^and_result26[140]^and_result26[141]^and_result26[142]^and_result26[143]^and_result26[144]^and_result26[145]^and_result26[146]^and_result26[147]^and_result26[148]^and_result26[149]^and_result26[150]^and_result26[151]^and_result26[152]^and_result26[153]^and_result26[154]^and_result26[155]^and_result26[156]^and_result26[157]^and_result26[158]^and_result26[159]^and_result26[160]^and_result26[161]^and_result26[162]^and_result26[163]^and_result26[164]^and_result26[165]^and_result26[166]^and_result26[167]^and_result26[168]^and_result26[169]^and_result26[170]^and_result26[171]^and_result26[172]^and_result26[173]^and_result26[174]^and_result26[175]^and_result26[176]^and_result26[177]^and_result26[178]^and_result26[179]^and_result26[180]^and_result26[181]^and_result26[182]^and_result26[183]^and_result26[184]^and_result26[185]^and_result26[186]^and_result26[187]^and_result26[188]^and_result26[189]^and_result26[190]^and_result26[191]^and_result26[192]^and_result26[193]^and_result26[194]^and_result26[195]^and_result26[196]^and_result26[197]^and_result26[198]^and_result26[199]^and_result26[200]^and_result26[201]^and_result26[202]^and_result26[203]^and_result26[204]^and_result26[205]^and_result26[206]^and_result26[207]^and_result26[208]^and_result26[209]^and_result26[210]^and_result26[211]^and_result26[212]^and_result26[213]^and_result26[214]^and_result26[215]^and_result26[216]^and_result26[217]^and_result26[218]^and_result26[219]^and_result26[220]^and_result26[221]^and_result26[222]^and_result26[223]^and_result26[224]^and_result26[225]^and_result26[226]^and_result26[227]^and_result26[228]^and_result26[229]^and_result26[230]^and_result26[231]^and_result26[232]^and_result26[233]^and_result26[234]^and_result26[235]^and_result26[236]^and_result26[237]^and_result26[238]^and_result26[239]^and_result26[240]^and_result26[241]^and_result26[242]^and_result26[243]^and_result26[244]^and_result26[245]^and_result26[246]^and_result26[247]^and_result26[248]^and_result26[249]^and_result26[250]^and_result26[251]^and_result26[252]^and_result26[253]^and_result26[254];
assign key[27]=and_result27[0]^and_result27[1]^and_result27[2]^and_result27[3]^and_result27[4]^and_result27[5]^and_result27[6]^and_result27[7]^and_result27[8]^and_result27[9]^and_result27[10]^and_result27[11]^and_result27[12]^and_result27[13]^and_result27[14]^and_result27[15]^and_result27[16]^and_result27[17]^and_result27[18]^and_result27[19]^and_result27[20]^and_result27[21]^and_result27[22]^and_result27[23]^and_result27[24]^and_result27[25]^and_result27[26]^and_result27[27]^and_result27[28]^and_result27[29]^and_result27[30]^and_result27[31]^and_result27[32]^and_result27[33]^and_result27[34]^and_result27[35]^and_result27[36]^and_result27[37]^and_result27[38]^and_result27[39]^and_result27[40]^and_result27[41]^and_result27[42]^and_result27[43]^and_result27[44]^and_result27[45]^and_result27[46]^and_result27[47]^and_result27[48]^and_result27[49]^and_result27[50]^and_result27[51]^and_result27[52]^and_result27[53]^and_result27[54]^and_result27[55]^and_result27[56]^and_result27[57]^and_result27[58]^and_result27[59]^and_result27[60]^and_result27[61]^and_result27[62]^and_result27[63]^and_result27[64]^and_result27[65]^and_result27[66]^and_result27[67]^and_result27[68]^and_result27[69]^and_result27[70]^and_result27[71]^and_result27[72]^and_result27[73]^and_result27[74]^and_result27[75]^and_result27[76]^and_result27[77]^and_result27[78]^and_result27[79]^and_result27[80]^and_result27[81]^and_result27[82]^and_result27[83]^and_result27[84]^and_result27[85]^and_result27[86]^and_result27[87]^and_result27[88]^and_result27[89]^and_result27[90]^and_result27[91]^and_result27[92]^and_result27[93]^and_result27[94]^and_result27[95]^and_result27[96]^and_result27[97]^and_result27[98]^and_result27[99]^and_result27[100]^and_result27[101]^and_result27[102]^and_result27[103]^and_result27[104]^and_result27[105]^and_result27[106]^and_result27[107]^and_result27[108]^and_result27[109]^and_result27[110]^and_result27[111]^and_result27[112]^and_result27[113]^and_result27[114]^and_result27[115]^and_result27[116]^and_result27[117]^and_result27[118]^and_result27[119]^and_result27[120]^and_result27[121]^and_result27[122]^and_result27[123]^and_result27[124]^and_result27[125]^and_result27[126]^and_result27[127]^and_result27[128]^and_result27[129]^and_result27[130]^and_result27[131]^and_result27[132]^and_result27[133]^and_result27[134]^and_result27[135]^and_result27[136]^and_result27[137]^and_result27[138]^and_result27[139]^and_result27[140]^and_result27[141]^and_result27[142]^and_result27[143]^and_result27[144]^and_result27[145]^and_result27[146]^and_result27[147]^and_result27[148]^and_result27[149]^and_result27[150]^and_result27[151]^and_result27[152]^and_result27[153]^and_result27[154]^and_result27[155]^and_result27[156]^and_result27[157]^and_result27[158]^and_result27[159]^and_result27[160]^and_result27[161]^and_result27[162]^and_result27[163]^and_result27[164]^and_result27[165]^and_result27[166]^and_result27[167]^and_result27[168]^and_result27[169]^and_result27[170]^and_result27[171]^and_result27[172]^and_result27[173]^and_result27[174]^and_result27[175]^and_result27[176]^and_result27[177]^and_result27[178]^and_result27[179]^and_result27[180]^and_result27[181]^and_result27[182]^and_result27[183]^and_result27[184]^and_result27[185]^and_result27[186]^and_result27[187]^and_result27[188]^and_result27[189]^and_result27[190]^and_result27[191]^and_result27[192]^and_result27[193]^and_result27[194]^and_result27[195]^and_result27[196]^and_result27[197]^and_result27[198]^and_result27[199]^and_result27[200]^and_result27[201]^and_result27[202]^and_result27[203]^and_result27[204]^and_result27[205]^and_result27[206]^and_result27[207]^and_result27[208]^and_result27[209]^and_result27[210]^and_result27[211]^and_result27[212]^and_result27[213]^and_result27[214]^and_result27[215]^and_result27[216]^and_result27[217]^and_result27[218]^and_result27[219]^and_result27[220]^and_result27[221]^and_result27[222]^and_result27[223]^and_result27[224]^and_result27[225]^and_result27[226]^and_result27[227]^and_result27[228]^and_result27[229]^and_result27[230]^and_result27[231]^and_result27[232]^and_result27[233]^and_result27[234]^and_result27[235]^and_result27[236]^and_result27[237]^and_result27[238]^and_result27[239]^and_result27[240]^and_result27[241]^and_result27[242]^and_result27[243]^and_result27[244]^and_result27[245]^and_result27[246]^and_result27[247]^and_result27[248]^and_result27[249]^and_result27[250]^and_result27[251]^and_result27[252]^and_result27[253]^and_result27[254];
assign key[28]=and_result28[0]^and_result28[1]^and_result28[2]^and_result28[3]^and_result28[4]^and_result28[5]^and_result28[6]^and_result28[7]^and_result28[8]^and_result28[9]^and_result28[10]^and_result28[11]^and_result28[12]^and_result28[13]^and_result28[14]^and_result28[15]^and_result28[16]^and_result28[17]^and_result28[18]^and_result28[19]^and_result28[20]^and_result28[21]^and_result28[22]^and_result28[23]^and_result28[24]^and_result28[25]^and_result28[26]^and_result28[27]^and_result28[28]^and_result28[29]^and_result28[30]^and_result28[31]^and_result28[32]^and_result28[33]^and_result28[34]^and_result28[35]^and_result28[36]^and_result28[37]^and_result28[38]^and_result28[39]^and_result28[40]^and_result28[41]^and_result28[42]^and_result28[43]^and_result28[44]^and_result28[45]^and_result28[46]^and_result28[47]^and_result28[48]^and_result28[49]^and_result28[50]^and_result28[51]^and_result28[52]^and_result28[53]^and_result28[54]^and_result28[55]^and_result28[56]^and_result28[57]^and_result28[58]^and_result28[59]^and_result28[60]^and_result28[61]^and_result28[62]^and_result28[63]^and_result28[64]^and_result28[65]^and_result28[66]^and_result28[67]^and_result28[68]^and_result28[69]^and_result28[70]^and_result28[71]^and_result28[72]^and_result28[73]^and_result28[74]^and_result28[75]^and_result28[76]^and_result28[77]^and_result28[78]^and_result28[79]^and_result28[80]^and_result28[81]^and_result28[82]^and_result28[83]^and_result28[84]^and_result28[85]^and_result28[86]^and_result28[87]^and_result28[88]^and_result28[89]^and_result28[90]^and_result28[91]^and_result28[92]^and_result28[93]^and_result28[94]^and_result28[95]^and_result28[96]^and_result28[97]^and_result28[98]^and_result28[99]^and_result28[100]^and_result28[101]^and_result28[102]^and_result28[103]^and_result28[104]^and_result28[105]^and_result28[106]^and_result28[107]^and_result28[108]^and_result28[109]^and_result28[110]^and_result28[111]^and_result28[112]^and_result28[113]^and_result28[114]^and_result28[115]^and_result28[116]^and_result28[117]^and_result28[118]^and_result28[119]^and_result28[120]^and_result28[121]^and_result28[122]^and_result28[123]^and_result28[124]^and_result28[125]^and_result28[126]^and_result28[127]^and_result28[128]^and_result28[129]^and_result28[130]^and_result28[131]^and_result28[132]^and_result28[133]^and_result28[134]^and_result28[135]^and_result28[136]^and_result28[137]^and_result28[138]^and_result28[139]^and_result28[140]^and_result28[141]^and_result28[142]^and_result28[143]^and_result28[144]^and_result28[145]^and_result28[146]^and_result28[147]^and_result28[148]^and_result28[149]^and_result28[150]^and_result28[151]^and_result28[152]^and_result28[153]^and_result28[154]^and_result28[155]^and_result28[156]^and_result28[157]^and_result28[158]^and_result28[159]^and_result28[160]^and_result28[161]^and_result28[162]^and_result28[163]^and_result28[164]^and_result28[165]^and_result28[166]^and_result28[167]^and_result28[168]^and_result28[169]^and_result28[170]^and_result28[171]^and_result28[172]^and_result28[173]^and_result28[174]^and_result28[175]^and_result28[176]^and_result28[177]^and_result28[178]^and_result28[179]^and_result28[180]^and_result28[181]^and_result28[182]^and_result28[183]^and_result28[184]^and_result28[185]^and_result28[186]^and_result28[187]^and_result28[188]^and_result28[189]^and_result28[190]^and_result28[191]^and_result28[192]^and_result28[193]^and_result28[194]^and_result28[195]^and_result28[196]^and_result28[197]^and_result28[198]^and_result28[199]^and_result28[200]^and_result28[201]^and_result28[202]^and_result28[203]^and_result28[204]^and_result28[205]^and_result28[206]^and_result28[207]^and_result28[208]^and_result28[209]^and_result28[210]^and_result28[211]^and_result28[212]^and_result28[213]^and_result28[214]^and_result28[215]^and_result28[216]^and_result28[217]^and_result28[218]^and_result28[219]^and_result28[220]^and_result28[221]^and_result28[222]^and_result28[223]^and_result28[224]^and_result28[225]^and_result28[226]^and_result28[227]^and_result28[228]^and_result28[229]^and_result28[230]^and_result28[231]^and_result28[232]^and_result28[233]^and_result28[234]^and_result28[235]^and_result28[236]^and_result28[237]^and_result28[238]^and_result28[239]^and_result28[240]^and_result28[241]^and_result28[242]^and_result28[243]^and_result28[244]^and_result28[245]^and_result28[246]^and_result28[247]^and_result28[248]^and_result28[249]^and_result28[250]^and_result28[251]^and_result28[252]^and_result28[253]^and_result28[254];
assign key[29]=and_result29[0]^and_result29[1]^and_result29[2]^and_result29[3]^and_result29[4]^and_result29[5]^and_result29[6]^and_result29[7]^and_result29[8]^and_result29[9]^and_result29[10]^and_result29[11]^and_result29[12]^and_result29[13]^and_result29[14]^and_result29[15]^and_result29[16]^and_result29[17]^and_result29[18]^and_result29[19]^and_result29[20]^and_result29[21]^and_result29[22]^and_result29[23]^and_result29[24]^and_result29[25]^and_result29[26]^and_result29[27]^and_result29[28]^and_result29[29]^and_result29[30]^and_result29[31]^and_result29[32]^and_result29[33]^and_result29[34]^and_result29[35]^and_result29[36]^and_result29[37]^and_result29[38]^and_result29[39]^and_result29[40]^and_result29[41]^and_result29[42]^and_result29[43]^and_result29[44]^and_result29[45]^and_result29[46]^and_result29[47]^and_result29[48]^and_result29[49]^and_result29[50]^and_result29[51]^and_result29[52]^and_result29[53]^and_result29[54]^and_result29[55]^and_result29[56]^and_result29[57]^and_result29[58]^and_result29[59]^and_result29[60]^and_result29[61]^and_result29[62]^and_result29[63]^and_result29[64]^and_result29[65]^and_result29[66]^and_result29[67]^and_result29[68]^and_result29[69]^and_result29[70]^and_result29[71]^and_result29[72]^and_result29[73]^and_result29[74]^and_result29[75]^and_result29[76]^and_result29[77]^and_result29[78]^and_result29[79]^and_result29[80]^and_result29[81]^and_result29[82]^and_result29[83]^and_result29[84]^and_result29[85]^and_result29[86]^and_result29[87]^and_result29[88]^and_result29[89]^and_result29[90]^and_result29[91]^and_result29[92]^and_result29[93]^and_result29[94]^and_result29[95]^and_result29[96]^and_result29[97]^and_result29[98]^and_result29[99]^and_result29[100]^and_result29[101]^and_result29[102]^and_result29[103]^and_result29[104]^and_result29[105]^and_result29[106]^and_result29[107]^and_result29[108]^and_result29[109]^and_result29[110]^and_result29[111]^and_result29[112]^and_result29[113]^and_result29[114]^and_result29[115]^and_result29[116]^and_result29[117]^and_result29[118]^and_result29[119]^and_result29[120]^and_result29[121]^and_result29[122]^and_result29[123]^and_result29[124]^and_result29[125]^and_result29[126]^and_result29[127]^and_result29[128]^and_result29[129]^and_result29[130]^and_result29[131]^and_result29[132]^and_result29[133]^and_result29[134]^and_result29[135]^and_result29[136]^and_result29[137]^and_result29[138]^and_result29[139]^and_result29[140]^and_result29[141]^and_result29[142]^and_result29[143]^and_result29[144]^and_result29[145]^and_result29[146]^and_result29[147]^and_result29[148]^and_result29[149]^and_result29[150]^and_result29[151]^and_result29[152]^and_result29[153]^and_result29[154]^and_result29[155]^and_result29[156]^and_result29[157]^and_result29[158]^and_result29[159]^and_result29[160]^and_result29[161]^and_result29[162]^and_result29[163]^and_result29[164]^and_result29[165]^and_result29[166]^and_result29[167]^and_result29[168]^and_result29[169]^and_result29[170]^and_result29[171]^and_result29[172]^and_result29[173]^and_result29[174]^and_result29[175]^and_result29[176]^and_result29[177]^and_result29[178]^and_result29[179]^and_result29[180]^and_result29[181]^and_result29[182]^and_result29[183]^and_result29[184]^and_result29[185]^and_result29[186]^and_result29[187]^and_result29[188]^and_result29[189]^and_result29[190]^and_result29[191]^and_result29[192]^and_result29[193]^and_result29[194]^and_result29[195]^and_result29[196]^and_result29[197]^and_result29[198]^and_result29[199]^and_result29[200]^and_result29[201]^and_result29[202]^and_result29[203]^and_result29[204]^and_result29[205]^and_result29[206]^and_result29[207]^and_result29[208]^and_result29[209]^and_result29[210]^and_result29[211]^and_result29[212]^and_result29[213]^and_result29[214]^and_result29[215]^and_result29[216]^and_result29[217]^and_result29[218]^and_result29[219]^and_result29[220]^and_result29[221]^and_result29[222]^and_result29[223]^and_result29[224]^and_result29[225]^and_result29[226]^and_result29[227]^and_result29[228]^and_result29[229]^and_result29[230]^and_result29[231]^and_result29[232]^and_result29[233]^and_result29[234]^and_result29[235]^and_result29[236]^and_result29[237]^and_result29[238]^and_result29[239]^and_result29[240]^and_result29[241]^and_result29[242]^and_result29[243]^and_result29[244]^and_result29[245]^and_result29[246]^and_result29[247]^and_result29[248]^and_result29[249]^and_result29[250]^and_result29[251]^and_result29[252]^and_result29[253]^and_result29[254];
assign key[30]=and_result30[0]^and_result30[1]^and_result30[2]^and_result30[3]^and_result30[4]^and_result30[5]^and_result30[6]^and_result30[7]^and_result30[8]^and_result30[9]^and_result30[10]^and_result30[11]^and_result30[12]^and_result30[13]^and_result30[14]^and_result30[15]^and_result30[16]^and_result30[17]^and_result30[18]^and_result30[19]^and_result30[20]^and_result30[21]^and_result30[22]^and_result30[23]^and_result30[24]^and_result30[25]^and_result30[26]^and_result30[27]^and_result30[28]^and_result30[29]^and_result30[30]^and_result30[31]^and_result30[32]^and_result30[33]^and_result30[34]^and_result30[35]^and_result30[36]^and_result30[37]^and_result30[38]^and_result30[39]^and_result30[40]^and_result30[41]^and_result30[42]^and_result30[43]^and_result30[44]^and_result30[45]^and_result30[46]^and_result30[47]^and_result30[48]^and_result30[49]^and_result30[50]^and_result30[51]^and_result30[52]^and_result30[53]^and_result30[54]^and_result30[55]^and_result30[56]^and_result30[57]^and_result30[58]^and_result30[59]^and_result30[60]^and_result30[61]^and_result30[62]^and_result30[63]^and_result30[64]^and_result30[65]^and_result30[66]^and_result30[67]^and_result30[68]^and_result30[69]^and_result30[70]^and_result30[71]^and_result30[72]^and_result30[73]^and_result30[74]^and_result30[75]^and_result30[76]^and_result30[77]^and_result30[78]^and_result30[79]^and_result30[80]^and_result30[81]^and_result30[82]^and_result30[83]^and_result30[84]^and_result30[85]^and_result30[86]^and_result30[87]^and_result30[88]^and_result30[89]^and_result30[90]^and_result30[91]^and_result30[92]^and_result30[93]^and_result30[94]^and_result30[95]^and_result30[96]^and_result30[97]^and_result30[98]^and_result30[99]^and_result30[100]^and_result30[101]^and_result30[102]^and_result30[103]^and_result30[104]^and_result30[105]^and_result30[106]^and_result30[107]^and_result30[108]^and_result30[109]^and_result30[110]^and_result30[111]^and_result30[112]^and_result30[113]^and_result30[114]^and_result30[115]^and_result30[116]^and_result30[117]^and_result30[118]^and_result30[119]^and_result30[120]^and_result30[121]^and_result30[122]^and_result30[123]^and_result30[124]^and_result30[125]^and_result30[126]^and_result30[127]^and_result30[128]^and_result30[129]^and_result30[130]^and_result30[131]^and_result30[132]^and_result30[133]^and_result30[134]^and_result30[135]^and_result30[136]^and_result30[137]^and_result30[138]^and_result30[139]^and_result30[140]^and_result30[141]^and_result30[142]^and_result30[143]^and_result30[144]^and_result30[145]^and_result30[146]^and_result30[147]^and_result30[148]^and_result30[149]^and_result30[150]^and_result30[151]^and_result30[152]^and_result30[153]^and_result30[154]^and_result30[155]^and_result30[156]^and_result30[157]^and_result30[158]^and_result30[159]^and_result30[160]^and_result30[161]^and_result30[162]^and_result30[163]^and_result30[164]^and_result30[165]^and_result30[166]^and_result30[167]^and_result30[168]^and_result30[169]^and_result30[170]^and_result30[171]^and_result30[172]^and_result30[173]^and_result30[174]^and_result30[175]^and_result30[176]^and_result30[177]^and_result30[178]^and_result30[179]^and_result30[180]^and_result30[181]^and_result30[182]^and_result30[183]^and_result30[184]^and_result30[185]^and_result30[186]^and_result30[187]^and_result30[188]^and_result30[189]^and_result30[190]^and_result30[191]^and_result30[192]^and_result30[193]^and_result30[194]^and_result30[195]^and_result30[196]^and_result30[197]^and_result30[198]^and_result30[199]^and_result30[200]^and_result30[201]^and_result30[202]^and_result30[203]^and_result30[204]^and_result30[205]^and_result30[206]^and_result30[207]^and_result30[208]^and_result30[209]^and_result30[210]^and_result30[211]^and_result30[212]^and_result30[213]^and_result30[214]^and_result30[215]^and_result30[216]^and_result30[217]^and_result30[218]^and_result30[219]^and_result30[220]^and_result30[221]^and_result30[222]^and_result30[223]^and_result30[224]^and_result30[225]^and_result30[226]^and_result30[227]^and_result30[228]^and_result30[229]^and_result30[230]^and_result30[231]^and_result30[232]^and_result30[233]^and_result30[234]^and_result30[235]^and_result30[236]^and_result30[237]^and_result30[238]^and_result30[239]^and_result30[240]^and_result30[241]^and_result30[242]^and_result30[243]^and_result30[244]^and_result30[245]^and_result30[246]^and_result30[247]^and_result30[248]^and_result30[249]^and_result30[250]^and_result30[251]^and_result30[252]^and_result30[253]^and_result30[254];
assign key[31]=and_result31[0]^and_result31[1]^and_result31[2]^and_result31[3]^and_result31[4]^and_result31[5]^and_result31[6]^and_result31[7]^and_result31[8]^and_result31[9]^and_result31[10]^and_result31[11]^and_result31[12]^and_result31[13]^and_result31[14]^and_result31[15]^and_result31[16]^and_result31[17]^and_result31[18]^and_result31[19]^and_result31[20]^and_result31[21]^and_result31[22]^and_result31[23]^and_result31[24]^and_result31[25]^and_result31[26]^and_result31[27]^and_result31[28]^and_result31[29]^and_result31[30]^and_result31[31]^and_result31[32]^and_result31[33]^and_result31[34]^and_result31[35]^and_result31[36]^and_result31[37]^and_result31[38]^and_result31[39]^and_result31[40]^and_result31[41]^and_result31[42]^and_result31[43]^and_result31[44]^and_result31[45]^and_result31[46]^and_result31[47]^and_result31[48]^and_result31[49]^and_result31[50]^and_result31[51]^and_result31[52]^and_result31[53]^and_result31[54]^and_result31[55]^and_result31[56]^and_result31[57]^and_result31[58]^and_result31[59]^and_result31[60]^and_result31[61]^and_result31[62]^and_result31[63]^and_result31[64]^and_result31[65]^and_result31[66]^and_result31[67]^and_result31[68]^and_result31[69]^and_result31[70]^and_result31[71]^and_result31[72]^and_result31[73]^and_result31[74]^and_result31[75]^and_result31[76]^and_result31[77]^and_result31[78]^and_result31[79]^and_result31[80]^and_result31[81]^and_result31[82]^and_result31[83]^and_result31[84]^and_result31[85]^and_result31[86]^and_result31[87]^and_result31[88]^and_result31[89]^and_result31[90]^and_result31[91]^and_result31[92]^and_result31[93]^and_result31[94]^and_result31[95]^and_result31[96]^and_result31[97]^and_result31[98]^and_result31[99]^and_result31[100]^and_result31[101]^and_result31[102]^and_result31[103]^and_result31[104]^and_result31[105]^and_result31[106]^and_result31[107]^and_result31[108]^and_result31[109]^and_result31[110]^and_result31[111]^and_result31[112]^and_result31[113]^and_result31[114]^and_result31[115]^and_result31[116]^and_result31[117]^and_result31[118]^and_result31[119]^and_result31[120]^and_result31[121]^and_result31[122]^and_result31[123]^and_result31[124]^and_result31[125]^and_result31[126]^and_result31[127]^and_result31[128]^and_result31[129]^and_result31[130]^and_result31[131]^and_result31[132]^and_result31[133]^and_result31[134]^and_result31[135]^and_result31[136]^and_result31[137]^and_result31[138]^and_result31[139]^and_result31[140]^and_result31[141]^and_result31[142]^and_result31[143]^and_result31[144]^and_result31[145]^and_result31[146]^and_result31[147]^and_result31[148]^and_result31[149]^and_result31[150]^and_result31[151]^and_result31[152]^and_result31[153]^and_result31[154]^and_result31[155]^and_result31[156]^and_result31[157]^and_result31[158]^and_result31[159]^and_result31[160]^and_result31[161]^and_result31[162]^and_result31[163]^and_result31[164]^and_result31[165]^and_result31[166]^and_result31[167]^and_result31[168]^and_result31[169]^and_result31[170]^and_result31[171]^and_result31[172]^and_result31[173]^and_result31[174]^and_result31[175]^and_result31[176]^and_result31[177]^and_result31[178]^and_result31[179]^and_result31[180]^and_result31[181]^and_result31[182]^and_result31[183]^and_result31[184]^and_result31[185]^and_result31[186]^and_result31[187]^and_result31[188]^and_result31[189]^and_result31[190]^and_result31[191]^and_result31[192]^and_result31[193]^and_result31[194]^and_result31[195]^and_result31[196]^and_result31[197]^and_result31[198]^and_result31[199]^and_result31[200]^and_result31[201]^and_result31[202]^and_result31[203]^and_result31[204]^and_result31[205]^and_result31[206]^and_result31[207]^and_result31[208]^and_result31[209]^and_result31[210]^and_result31[211]^and_result31[212]^and_result31[213]^and_result31[214]^and_result31[215]^and_result31[216]^and_result31[217]^and_result31[218]^and_result31[219]^and_result31[220]^and_result31[221]^and_result31[222]^and_result31[223]^and_result31[224]^and_result31[225]^and_result31[226]^and_result31[227]^and_result31[228]^and_result31[229]^and_result31[230]^and_result31[231]^and_result31[232]^and_result31[233]^and_result31[234]^and_result31[235]^and_result31[236]^and_result31[237]^and_result31[238]^and_result31[239]^and_result31[240]^and_result31[241]^and_result31[242]^and_result31[243]^and_result31[244]^and_result31[245]^and_result31[246]^and_result31[247]^and_result31[248]^and_result31[249]^and_result31[250]^and_result31[251]^and_result31[252]^and_result31[253]^and_result31[254];
assign key[32]=and_result32[0]^and_result32[1]^and_result32[2]^and_result32[3]^and_result32[4]^and_result32[5]^and_result32[6]^and_result32[7]^and_result32[8]^and_result32[9]^and_result32[10]^and_result32[11]^and_result32[12]^and_result32[13]^and_result32[14]^and_result32[15]^and_result32[16]^and_result32[17]^and_result32[18]^and_result32[19]^and_result32[20]^and_result32[21]^and_result32[22]^and_result32[23]^and_result32[24]^and_result32[25]^and_result32[26]^and_result32[27]^and_result32[28]^and_result32[29]^and_result32[30]^and_result32[31]^and_result32[32]^and_result32[33]^and_result32[34]^and_result32[35]^and_result32[36]^and_result32[37]^and_result32[38]^and_result32[39]^and_result32[40]^and_result32[41]^and_result32[42]^and_result32[43]^and_result32[44]^and_result32[45]^and_result32[46]^and_result32[47]^and_result32[48]^and_result32[49]^and_result32[50]^and_result32[51]^and_result32[52]^and_result32[53]^and_result32[54]^and_result32[55]^and_result32[56]^and_result32[57]^and_result32[58]^and_result32[59]^and_result32[60]^and_result32[61]^and_result32[62]^and_result32[63]^and_result32[64]^and_result32[65]^and_result32[66]^and_result32[67]^and_result32[68]^and_result32[69]^and_result32[70]^and_result32[71]^and_result32[72]^and_result32[73]^and_result32[74]^and_result32[75]^and_result32[76]^and_result32[77]^and_result32[78]^and_result32[79]^and_result32[80]^and_result32[81]^and_result32[82]^and_result32[83]^and_result32[84]^and_result32[85]^and_result32[86]^and_result32[87]^and_result32[88]^and_result32[89]^and_result32[90]^and_result32[91]^and_result32[92]^and_result32[93]^and_result32[94]^and_result32[95]^and_result32[96]^and_result32[97]^and_result32[98]^and_result32[99]^and_result32[100]^and_result32[101]^and_result32[102]^and_result32[103]^and_result32[104]^and_result32[105]^and_result32[106]^and_result32[107]^and_result32[108]^and_result32[109]^and_result32[110]^and_result32[111]^and_result32[112]^and_result32[113]^and_result32[114]^and_result32[115]^and_result32[116]^and_result32[117]^and_result32[118]^and_result32[119]^and_result32[120]^and_result32[121]^and_result32[122]^and_result32[123]^and_result32[124]^and_result32[125]^and_result32[126]^and_result32[127]^and_result32[128]^and_result32[129]^and_result32[130]^and_result32[131]^and_result32[132]^and_result32[133]^and_result32[134]^and_result32[135]^and_result32[136]^and_result32[137]^and_result32[138]^and_result32[139]^and_result32[140]^and_result32[141]^and_result32[142]^and_result32[143]^and_result32[144]^and_result32[145]^and_result32[146]^and_result32[147]^and_result32[148]^and_result32[149]^and_result32[150]^and_result32[151]^and_result32[152]^and_result32[153]^and_result32[154]^and_result32[155]^and_result32[156]^and_result32[157]^and_result32[158]^and_result32[159]^and_result32[160]^and_result32[161]^and_result32[162]^and_result32[163]^and_result32[164]^and_result32[165]^and_result32[166]^and_result32[167]^and_result32[168]^and_result32[169]^and_result32[170]^and_result32[171]^and_result32[172]^and_result32[173]^and_result32[174]^and_result32[175]^and_result32[176]^and_result32[177]^and_result32[178]^and_result32[179]^and_result32[180]^and_result32[181]^and_result32[182]^and_result32[183]^and_result32[184]^and_result32[185]^and_result32[186]^and_result32[187]^and_result32[188]^and_result32[189]^and_result32[190]^and_result32[191]^and_result32[192]^and_result32[193]^and_result32[194]^and_result32[195]^and_result32[196]^and_result32[197]^and_result32[198]^and_result32[199]^and_result32[200]^and_result32[201]^and_result32[202]^and_result32[203]^and_result32[204]^and_result32[205]^and_result32[206]^and_result32[207]^and_result32[208]^and_result32[209]^and_result32[210]^and_result32[211]^and_result32[212]^and_result32[213]^and_result32[214]^and_result32[215]^and_result32[216]^and_result32[217]^and_result32[218]^and_result32[219]^and_result32[220]^and_result32[221]^and_result32[222]^and_result32[223]^and_result32[224]^and_result32[225]^and_result32[226]^and_result32[227]^and_result32[228]^and_result32[229]^and_result32[230]^and_result32[231]^and_result32[232]^and_result32[233]^and_result32[234]^and_result32[235]^and_result32[236]^and_result32[237]^and_result32[238]^and_result32[239]^and_result32[240]^and_result32[241]^and_result32[242]^and_result32[243]^and_result32[244]^and_result32[245]^and_result32[246]^and_result32[247]^and_result32[248]^and_result32[249]^and_result32[250]^and_result32[251]^and_result32[252]^and_result32[253]^and_result32[254];
assign key[33]=and_result33[0]^and_result33[1]^and_result33[2]^and_result33[3]^and_result33[4]^and_result33[5]^and_result33[6]^and_result33[7]^and_result33[8]^and_result33[9]^and_result33[10]^and_result33[11]^and_result33[12]^and_result33[13]^and_result33[14]^and_result33[15]^and_result33[16]^and_result33[17]^and_result33[18]^and_result33[19]^and_result33[20]^and_result33[21]^and_result33[22]^and_result33[23]^and_result33[24]^and_result33[25]^and_result33[26]^and_result33[27]^and_result33[28]^and_result33[29]^and_result33[30]^and_result33[31]^and_result33[32]^and_result33[33]^and_result33[34]^and_result33[35]^and_result33[36]^and_result33[37]^and_result33[38]^and_result33[39]^and_result33[40]^and_result33[41]^and_result33[42]^and_result33[43]^and_result33[44]^and_result33[45]^and_result33[46]^and_result33[47]^and_result33[48]^and_result33[49]^and_result33[50]^and_result33[51]^and_result33[52]^and_result33[53]^and_result33[54]^and_result33[55]^and_result33[56]^and_result33[57]^and_result33[58]^and_result33[59]^and_result33[60]^and_result33[61]^and_result33[62]^and_result33[63]^and_result33[64]^and_result33[65]^and_result33[66]^and_result33[67]^and_result33[68]^and_result33[69]^and_result33[70]^and_result33[71]^and_result33[72]^and_result33[73]^and_result33[74]^and_result33[75]^and_result33[76]^and_result33[77]^and_result33[78]^and_result33[79]^and_result33[80]^and_result33[81]^and_result33[82]^and_result33[83]^and_result33[84]^and_result33[85]^and_result33[86]^and_result33[87]^and_result33[88]^and_result33[89]^and_result33[90]^and_result33[91]^and_result33[92]^and_result33[93]^and_result33[94]^and_result33[95]^and_result33[96]^and_result33[97]^and_result33[98]^and_result33[99]^and_result33[100]^and_result33[101]^and_result33[102]^and_result33[103]^and_result33[104]^and_result33[105]^and_result33[106]^and_result33[107]^and_result33[108]^and_result33[109]^and_result33[110]^and_result33[111]^and_result33[112]^and_result33[113]^and_result33[114]^and_result33[115]^and_result33[116]^and_result33[117]^and_result33[118]^and_result33[119]^and_result33[120]^and_result33[121]^and_result33[122]^and_result33[123]^and_result33[124]^and_result33[125]^and_result33[126]^and_result33[127]^and_result33[128]^and_result33[129]^and_result33[130]^and_result33[131]^and_result33[132]^and_result33[133]^and_result33[134]^and_result33[135]^and_result33[136]^and_result33[137]^and_result33[138]^and_result33[139]^and_result33[140]^and_result33[141]^and_result33[142]^and_result33[143]^and_result33[144]^and_result33[145]^and_result33[146]^and_result33[147]^and_result33[148]^and_result33[149]^and_result33[150]^and_result33[151]^and_result33[152]^and_result33[153]^and_result33[154]^and_result33[155]^and_result33[156]^and_result33[157]^and_result33[158]^and_result33[159]^and_result33[160]^and_result33[161]^and_result33[162]^and_result33[163]^and_result33[164]^and_result33[165]^and_result33[166]^and_result33[167]^and_result33[168]^and_result33[169]^and_result33[170]^and_result33[171]^and_result33[172]^and_result33[173]^and_result33[174]^and_result33[175]^and_result33[176]^and_result33[177]^and_result33[178]^and_result33[179]^and_result33[180]^and_result33[181]^and_result33[182]^and_result33[183]^and_result33[184]^and_result33[185]^and_result33[186]^and_result33[187]^and_result33[188]^and_result33[189]^and_result33[190]^and_result33[191]^and_result33[192]^and_result33[193]^and_result33[194]^and_result33[195]^and_result33[196]^and_result33[197]^and_result33[198]^and_result33[199]^and_result33[200]^and_result33[201]^and_result33[202]^and_result33[203]^and_result33[204]^and_result33[205]^and_result33[206]^and_result33[207]^and_result33[208]^and_result33[209]^and_result33[210]^and_result33[211]^and_result33[212]^and_result33[213]^and_result33[214]^and_result33[215]^and_result33[216]^and_result33[217]^and_result33[218]^and_result33[219]^and_result33[220]^and_result33[221]^and_result33[222]^and_result33[223]^and_result33[224]^and_result33[225]^and_result33[226]^and_result33[227]^and_result33[228]^and_result33[229]^and_result33[230]^and_result33[231]^and_result33[232]^and_result33[233]^and_result33[234]^and_result33[235]^and_result33[236]^and_result33[237]^and_result33[238]^and_result33[239]^and_result33[240]^and_result33[241]^and_result33[242]^and_result33[243]^and_result33[244]^and_result33[245]^and_result33[246]^and_result33[247]^and_result33[248]^and_result33[249]^and_result33[250]^and_result33[251]^and_result33[252]^and_result33[253]^and_result33[254];
assign key[34]=and_result34[0]^and_result34[1]^and_result34[2]^and_result34[3]^and_result34[4]^and_result34[5]^and_result34[6]^and_result34[7]^and_result34[8]^and_result34[9]^and_result34[10]^and_result34[11]^and_result34[12]^and_result34[13]^and_result34[14]^and_result34[15]^and_result34[16]^and_result34[17]^and_result34[18]^and_result34[19]^and_result34[20]^and_result34[21]^and_result34[22]^and_result34[23]^and_result34[24]^and_result34[25]^and_result34[26]^and_result34[27]^and_result34[28]^and_result34[29]^and_result34[30]^and_result34[31]^and_result34[32]^and_result34[33]^and_result34[34]^and_result34[35]^and_result34[36]^and_result34[37]^and_result34[38]^and_result34[39]^and_result34[40]^and_result34[41]^and_result34[42]^and_result34[43]^and_result34[44]^and_result34[45]^and_result34[46]^and_result34[47]^and_result34[48]^and_result34[49]^and_result34[50]^and_result34[51]^and_result34[52]^and_result34[53]^and_result34[54]^and_result34[55]^and_result34[56]^and_result34[57]^and_result34[58]^and_result34[59]^and_result34[60]^and_result34[61]^and_result34[62]^and_result34[63]^and_result34[64]^and_result34[65]^and_result34[66]^and_result34[67]^and_result34[68]^and_result34[69]^and_result34[70]^and_result34[71]^and_result34[72]^and_result34[73]^and_result34[74]^and_result34[75]^and_result34[76]^and_result34[77]^and_result34[78]^and_result34[79]^and_result34[80]^and_result34[81]^and_result34[82]^and_result34[83]^and_result34[84]^and_result34[85]^and_result34[86]^and_result34[87]^and_result34[88]^and_result34[89]^and_result34[90]^and_result34[91]^and_result34[92]^and_result34[93]^and_result34[94]^and_result34[95]^and_result34[96]^and_result34[97]^and_result34[98]^and_result34[99]^and_result34[100]^and_result34[101]^and_result34[102]^and_result34[103]^and_result34[104]^and_result34[105]^and_result34[106]^and_result34[107]^and_result34[108]^and_result34[109]^and_result34[110]^and_result34[111]^and_result34[112]^and_result34[113]^and_result34[114]^and_result34[115]^and_result34[116]^and_result34[117]^and_result34[118]^and_result34[119]^and_result34[120]^and_result34[121]^and_result34[122]^and_result34[123]^and_result34[124]^and_result34[125]^and_result34[126]^and_result34[127]^and_result34[128]^and_result34[129]^and_result34[130]^and_result34[131]^and_result34[132]^and_result34[133]^and_result34[134]^and_result34[135]^and_result34[136]^and_result34[137]^and_result34[138]^and_result34[139]^and_result34[140]^and_result34[141]^and_result34[142]^and_result34[143]^and_result34[144]^and_result34[145]^and_result34[146]^and_result34[147]^and_result34[148]^and_result34[149]^and_result34[150]^and_result34[151]^and_result34[152]^and_result34[153]^and_result34[154]^and_result34[155]^and_result34[156]^and_result34[157]^and_result34[158]^and_result34[159]^and_result34[160]^and_result34[161]^and_result34[162]^and_result34[163]^and_result34[164]^and_result34[165]^and_result34[166]^and_result34[167]^and_result34[168]^and_result34[169]^and_result34[170]^and_result34[171]^and_result34[172]^and_result34[173]^and_result34[174]^and_result34[175]^and_result34[176]^and_result34[177]^and_result34[178]^and_result34[179]^and_result34[180]^and_result34[181]^and_result34[182]^and_result34[183]^and_result34[184]^and_result34[185]^and_result34[186]^and_result34[187]^and_result34[188]^and_result34[189]^and_result34[190]^and_result34[191]^and_result34[192]^and_result34[193]^and_result34[194]^and_result34[195]^and_result34[196]^and_result34[197]^and_result34[198]^and_result34[199]^and_result34[200]^and_result34[201]^and_result34[202]^and_result34[203]^and_result34[204]^and_result34[205]^and_result34[206]^and_result34[207]^and_result34[208]^and_result34[209]^and_result34[210]^and_result34[211]^and_result34[212]^and_result34[213]^and_result34[214]^and_result34[215]^and_result34[216]^and_result34[217]^and_result34[218]^and_result34[219]^and_result34[220]^and_result34[221]^and_result34[222]^and_result34[223]^and_result34[224]^and_result34[225]^and_result34[226]^and_result34[227]^and_result34[228]^and_result34[229]^and_result34[230]^and_result34[231]^and_result34[232]^and_result34[233]^and_result34[234]^and_result34[235]^and_result34[236]^and_result34[237]^and_result34[238]^and_result34[239]^and_result34[240]^and_result34[241]^and_result34[242]^and_result34[243]^and_result34[244]^and_result34[245]^and_result34[246]^and_result34[247]^and_result34[248]^and_result34[249]^and_result34[250]^and_result34[251]^and_result34[252]^and_result34[253]^and_result34[254];
assign key[35]=and_result35[0]^and_result35[1]^and_result35[2]^and_result35[3]^and_result35[4]^and_result35[5]^and_result35[6]^and_result35[7]^and_result35[8]^and_result35[9]^and_result35[10]^and_result35[11]^and_result35[12]^and_result35[13]^and_result35[14]^and_result35[15]^and_result35[16]^and_result35[17]^and_result35[18]^and_result35[19]^and_result35[20]^and_result35[21]^and_result35[22]^and_result35[23]^and_result35[24]^and_result35[25]^and_result35[26]^and_result35[27]^and_result35[28]^and_result35[29]^and_result35[30]^and_result35[31]^and_result35[32]^and_result35[33]^and_result35[34]^and_result35[35]^and_result35[36]^and_result35[37]^and_result35[38]^and_result35[39]^and_result35[40]^and_result35[41]^and_result35[42]^and_result35[43]^and_result35[44]^and_result35[45]^and_result35[46]^and_result35[47]^and_result35[48]^and_result35[49]^and_result35[50]^and_result35[51]^and_result35[52]^and_result35[53]^and_result35[54]^and_result35[55]^and_result35[56]^and_result35[57]^and_result35[58]^and_result35[59]^and_result35[60]^and_result35[61]^and_result35[62]^and_result35[63]^and_result35[64]^and_result35[65]^and_result35[66]^and_result35[67]^and_result35[68]^and_result35[69]^and_result35[70]^and_result35[71]^and_result35[72]^and_result35[73]^and_result35[74]^and_result35[75]^and_result35[76]^and_result35[77]^and_result35[78]^and_result35[79]^and_result35[80]^and_result35[81]^and_result35[82]^and_result35[83]^and_result35[84]^and_result35[85]^and_result35[86]^and_result35[87]^and_result35[88]^and_result35[89]^and_result35[90]^and_result35[91]^and_result35[92]^and_result35[93]^and_result35[94]^and_result35[95]^and_result35[96]^and_result35[97]^and_result35[98]^and_result35[99]^and_result35[100]^and_result35[101]^and_result35[102]^and_result35[103]^and_result35[104]^and_result35[105]^and_result35[106]^and_result35[107]^and_result35[108]^and_result35[109]^and_result35[110]^and_result35[111]^and_result35[112]^and_result35[113]^and_result35[114]^and_result35[115]^and_result35[116]^and_result35[117]^and_result35[118]^and_result35[119]^and_result35[120]^and_result35[121]^and_result35[122]^and_result35[123]^and_result35[124]^and_result35[125]^and_result35[126]^and_result35[127]^and_result35[128]^and_result35[129]^and_result35[130]^and_result35[131]^and_result35[132]^and_result35[133]^and_result35[134]^and_result35[135]^and_result35[136]^and_result35[137]^and_result35[138]^and_result35[139]^and_result35[140]^and_result35[141]^and_result35[142]^and_result35[143]^and_result35[144]^and_result35[145]^and_result35[146]^and_result35[147]^and_result35[148]^and_result35[149]^and_result35[150]^and_result35[151]^and_result35[152]^and_result35[153]^and_result35[154]^and_result35[155]^and_result35[156]^and_result35[157]^and_result35[158]^and_result35[159]^and_result35[160]^and_result35[161]^and_result35[162]^and_result35[163]^and_result35[164]^and_result35[165]^and_result35[166]^and_result35[167]^and_result35[168]^and_result35[169]^and_result35[170]^and_result35[171]^and_result35[172]^and_result35[173]^and_result35[174]^and_result35[175]^and_result35[176]^and_result35[177]^and_result35[178]^and_result35[179]^and_result35[180]^and_result35[181]^and_result35[182]^and_result35[183]^and_result35[184]^and_result35[185]^and_result35[186]^and_result35[187]^and_result35[188]^and_result35[189]^and_result35[190]^and_result35[191]^and_result35[192]^and_result35[193]^and_result35[194]^and_result35[195]^and_result35[196]^and_result35[197]^and_result35[198]^and_result35[199]^and_result35[200]^and_result35[201]^and_result35[202]^and_result35[203]^and_result35[204]^and_result35[205]^and_result35[206]^and_result35[207]^and_result35[208]^and_result35[209]^and_result35[210]^and_result35[211]^and_result35[212]^and_result35[213]^and_result35[214]^and_result35[215]^and_result35[216]^and_result35[217]^and_result35[218]^and_result35[219]^and_result35[220]^and_result35[221]^and_result35[222]^and_result35[223]^and_result35[224]^and_result35[225]^and_result35[226]^and_result35[227]^and_result35[228]^and_result35[229]^and_result35[230]^and_result35[231]^and_result35[232]^and_result35[233]^and_result35[234]^and_result35[235]^and_result35[236]^and_result35[237]^and_result35[238]^and_result35[239]^and_result35[240]^and_result35[241]^and_result35[242]^and_result35[243]^and_result35[244]^and_result35[245]^and_result35[246]^and_result35[247]^and_result35[248]^and_result35[249]^and_result35[250]^and_result35[251]^and_result35[252]^and_result35[253]^and_result35[254];
assign key[36]=and_result36[0]^and_result36[1]^and_result36[2]^and_result36[3]^and_result36[4]^and_result36[5]^and_result36[6]^and_result36[7]^and_result36[8]^and_result36[9]^and_result36[10]^and_result36[11]^and_result36[12]^and_result36[13]^and_result36[14]^and_result36[15]^and_result36[16]^and_result36[17]^and_result36[18]^and_result36[19]^and_result36[20]^and_result36[21]^and_result36[22]^and_result36[23]^and_result36[24]^and_result36[25]^and_result36[26]^and_result36[27]^and_result36[28]^and_result36[29]^and_result36[30]^and_result36[31]^and_result36[32]^and_result36[33]^and_result36[34]^and_result36[35]^and_result36[36]^and_result36[37]^and_result36[38]^and_result36[39]^and_result36[40]^and_result36[41]^and_result36[42]^and_result36[43]^and_result36[44]^and_result36[45]^and_result36[46]^and_result36[47]^and_result36[48]^and_result36[49]^and_result36[50]^and_result36[51]^and_result36[52]^and_result36[53]^and_result36[54]^and_result36[55]^and_result36[56]^and_result36[57]^and_result36[58]^and_result36[59]^and_result36[60]^and_result36[61]^and_result36[62]^and_result36[63]^and_result36[64]^and_result36[65]^and_result36[66]^and_result36[67]^and_result36[68]^and_result36[69]^and_result36[70]^and_result36[71]^and_result36[72]^and_result36[73]^and_result36[74]^and_result36[75]^and_result36[76]^and_result36[77]^and_result36[78]^and_result36[79]^and_result36[80]^and_result36[81]^and_result36[82]^and_result36[83]^and_result36[84]^and_result36[85]^and_result36[86]^and_result36[87]^and_result36[88]^and_result36[89]^and_result36[90]^and_result36[91]^and_result36[92]^and_result36[93]^and_result36[94]^and_result36[95]^and_result36[96]^and_result36[97]^and_result36[98]^and_result36[99]^and_result36[100]^and_result36[101]^and_result36[102]^and_result36[103]^and_result36[104]^and_result36[105]^and_result36[106]^and_result36[107]^and_result36[108]^and_result36[109]^and_result36[110]^and_result36[111]^and_result36[112]^and_result36[113]^and_result36[114]^and_result36[115]^and_result36[116]^and_result36[117]^and_result36[118]^and_result36[119]^and_result36[120]^and_result36[121]^and_result36[122]^and_result36[123]^and_result36[124]^and_result36[125]^and_result36[126]^and_result36[127]^and_result36[128]^and_result36[129]^and_result36[130]^and_result36[131]^and_result36[132]^and_result36[133]^and_result36[134]^and_result36[135]^and_result36[136]^and_result36[137]^and_result36[138]^and_result36[139]^and_result36[140]^and_result36[141]^and_result36[142]^and_result36[143]^and_result36[144]^and_result36[145]^and_result36[146]^and_result36[147]^and_result36[148]^and_result36[149]^and_result36[150]^and_result36[151]^and_result36[152]^and_result36[153]^and_result36[154]^and_result36[155]^and_result36[156]^and_result36[157]^and_result36[158]^and_result36[159]^and_result36[160]^and_result36[161]^and_result36[162]^and_result36[163]^and_result36[164]^and_result36[165]^and_result36[166]^and_result36[167]^and_result36[168]^and_result36[169]^and_result36[170]^and_result36[171]^and_result36[172]^and_result36[173]^and_result36[174]^and_result36[175]^and_result36[176]^and_result36[177]^and_result36[178]^and_result36[179]^and_result36[180]^and_result36[181]^and_result36[182]^and_result36[183]^and_result36[184]^and_result36[185]^and_result36[186]^and_result36[187]^and_result36[188]^and_result36[189]^and_result36[190]^and_result36[191]^and_result36[192]^and_result36[193]^and_result36[194]^and_result36[195]^and_result36[196]^and_result36[197]^and_result36[198]^and_result36[199]^and_result36[200]^and_result36[201]^and_result36[202]^and_result36[203]^and_result36[204]^and_result36[205]^and_result36[206]^and_result36[207]^and_result36[208]^and_result36[209]^and_result36[210]^and_result36[211]^and_result36[212]^and_result36[213]^and_result36[214]^and_result36[215]^and_result36[216]^and_result36[217]^and_result36[218]^and_result36[219]^and_result36[220]^and_result36[221]^and_result36[222]^and_result36[223]^and_result36[224]^and_result36[225]^and_result36[226]^and_result36[227]^and_result36[228]^and_result36[229]^and_result36[230]^and_result36[231]^and_result36[232]^and_result36[233]^and_result36[234]^and_result36[235]^and_result36[236]^and_result36[237]^and_result36[238]^and_result36[239]^and_result36[240]^and_result36[241]^and_result36[242]^and_result36[243]^and_result36[244]^and_result36[245]^and_result36[246]^and_result36[247]^and_result36[248]^and_result36[249]^and_result36[250]^and_result36[251]^and_result36[252]^and_result36[253]^and_result36[254];
assign key[37]=and_result37[0]^and_result37[1]^and_result37[2]^and_result37[3]^and_result37[4]^and_result37[5]^and_result37[6]^and_result37[7]^and_result37[8]^and_result37[9]^and_result37[10]^and_result37[11]^and_result37[12]^and_result37[13]^and_result37[14]^and_result37[15]^and_result37[16]^and_result37[17]^and_result37[18]^and_result37[19]^and_result37[20]^and_result37[21]^and_result37[22]^and_result37[23]^and_result37[24]^and_result37[25]^and_result37[26]^and_result37[27]^and_result37[28]^and_result37[29]^and_result37[30]^and_result37[31]^and_result37[32]^and_result37[33]^and_result37[34]^and_result37[35]^and_result37[36]^and_result37[37]^and_result37[38]^and_result37[39]^and_result37[40]^and_result37[41]^and_result37[42]^and_result37[43]^and_result37[44]^and_result37[45]^and_result37[46]^and_result37[47]^and_result37[48]^and_result37[49]^and_result37[50]^and_result37[51]^and_result37[52]^and_result37[53]^and_result37[54]^and_result37[55]^and_result37[56]^and_result37[57]^and_result37[58]^and_result37[59]^and_result37[60]^and_result37[61]^and_result37[62]^and_result37[63]^and_result37[64]^and_result37[65]^and_result37[66]^and_result37[67]^and_result37[68]^and_result37[69]^and_result37[70]^and_result37[71]^and_result37[72]^and_result37[73]^and_result37[74]^and_result37[75]^and_result37[76]^and_result37[77]^and_result37[78]^and_result37[79]^and_result37[80]^and_result37[81]^and_result37[82]^and_result37[83]^and_result37[84]^and_result37[85]^and_result37[86]^and_result37[87]^and_result37[88]^and_result37[89]^and_result37[90]^and_result37[91]^and_result37[92]^and_result37[93]^and_result37[94]^and_result37[95]^and_result37[96]^and_result37[97]^and_result37[98]^and_result37[99]^and_result37[100]^and_result37[101]^and_result37[102]^and_result37[103]^and_result37[104]^and_result37[105]^and_result37[106]^and_result37[107]^and_result37[108]^and_result37[109]^and_result37[110]^and_result37[111]^and_result37[112]^and_result37[113]^and_result37[114]^and_result37[115]^and_result37[116]^and_result37[117]^and_result37[118]^and_result37[119]^and_result37[120]^and_result37[121]^and_result37[122]^and_result37[123]^and_result37[124]^and_result37[125]^and_result37[126]^and_result37[127]^and_result37[128]^and_result37[129]^and_result37[130]^and_result37[131]^and_result37[132]^and_result37[133]^and_result37[134]^and_result37[135]^and_result37[136]^and_result37[137]^and_result37[138]^and_result37[139]^and_result37[140]^and_result37[141]^and_result37[142]^and_result37[143]^and_result37[144]^and_result37[145]^and_result37[146]^and_result37[147]^and_result37[148]^and_result37[149]^and_result37[150]^and_result37[151]^and_result37[152]^and_result37[153]^and_result37[154]^and_result37[155]^and_result37[156]^and_result37[157]^and_result37[158]^and_result37[159]^and_result37[160]^and_result37[161]^and_result37[162]^and_result37[163]^and_result37[164]^and_result37[165]^and_result37[166]^and_result37[167]^and_result37[168]^and_result37[169]^and_result37[170]^and_result37[171]^and_result37[172]^and_result37[173]^and_result37[174]^and_result37[175]^and_result37[176]^and_result37[177]^and_result37[178]^and_result37[179]^and_result37[180]^and_result37[181]^and_result37[182]^and_result37[183]^and_result37[184]^and_result37[185]^and_result37[186]^and_result37[187]^and_result37[188]^and_result37[189]^and_result37[190]^and_result37[191]^and_result37[192]^and_result37[193]^and_result37[194]^and_result37[195]^and_result37[196]^and_result37[197]^and_result37[198]^and_result37[199]^and_result37[200]^and_result37[201]^and_result37[202]^and_result37[203]^and_result37[204]^and_result37[205]^and_result37[206]^and_result37[207]^and_result37[208]^and_result37[209]^and_result37[210]^and_result37[211]^and_result37[212]^and_result37[213]^and_result37[214]^and_result37[215]^and_result37[216]^and_result37[217]^and_result37[218]^and_result37[219]^and_result37[220]^and_result37[221]^and_result37[222]^and_result37[223]^and_result37[224]^and_result37[225]^and_result37[226]^and_result37[227]^and_result37[228]^and_result37[229]^and_result37[230]^and_result37[231]^and_result37[232]^and_result37[233]^and_result37[234]^and_result37[235]^and_result37[236]^and_result37[237]^and_result37[238]^and_result37[239]^and_result37[240]^and_result37[241]^and_result37[242]^and_result37[243]^and_result37[244]^and_result37[245]^and_result37[246]^and_result37[247]^and_result37[248]^and_result37[249]^and_result37[250]^and_result37[251]^and_result37[252]^and_result37[253]^and_result37[254];
assign key[38]=and_result38[0]^and_result38[1]^and_result38[2]^and_result38[3]^and_result38[4]^and_result38[5]^and_result38[6]^and_result38[7]^and_result38[8]^and_result38[9]^and_result38[10]^and_result38[11]^and_result38[12]^and_result38[13]^and_result38[14]^and_result38[15]^and_result38[16]^and_result38[17]^and_result38[18]^and_result38[19]^and_result38[20]^and_result38[21]^and_result38[22]^and_result38[23]^and_result38[24]^and_result38[25]^and_result38[26]^and_result38[27]^and_result38[28]^and_result38[29]^and_result38[30]^and_result38[31]^and_result38[32]^and_result38[33]^and_result38[34]^and_result38[35]^and_result38[36]^and_result38[37]^and_result38[38]^and_result38[39]^and_result38[40]^and_result38[41]^and_result38[42]^and_result38[43]^and_result38[44]^and_result38[45]^and_result38[46]^and_result38[47]^and_result38[48]^and_result38[49]^and_result38[50]^and_result38[51]^and_result38[52]^and_result38[53]^and_result38[54]^and_result38[55]^and_result38[56]^and_result38[57]^and_result38[58]^and_result38[59]^and_result38[60]^and_result38[61]^and_result38[62]^and_result38[63]^and_result38[64]^and_result38[65]^and_result38[66]^and_result38[67]^and_result38[68]^and_result38[69]^and_result38[70]^and_result38[71]^and_result38[72]^and_result38[73]^and_result38[74]^and_result38[75]^and_result38[76]^and_result38[77]^and_result38[78]^and_result38[79]^and_result38[80]^and_result38[81]^and_result38[82]^and_result38[83]^and_result38[84]^and_result38[85]^and_result38[86]^and_result38[87]^and_result38[88]^and_result38[89]^and_result38[90]^and_result38[91]^and_result38[92]^and_result38[93]^and_result38[94]^and_result38[95]^and_result38[96]^and_result38[97]^and_result38[98]^and_result38[99]^and_result38[100]^and_result38[101]^and_result38[102]^and_result38[103]^and_result38[104]^and_result38[105]^and_result38[106]^and_result38[107]^and_result38[108]^and_result38[109]^and_result38[110]^and_result38[111]^and_result38[112]^and_result38[113]^and_result38[114]^and_result38[115]^and_result38[116]^and_result38[117]^and_result38[118]^and_result38[119]^and_result38[120]^and_result38[121]^and_result38[122]^and_result38[123]^and_result38[124]^and_result38[125]^and_result38[126]^and_result38[127]^and_result38[128]^and_result38[129]^and_result38[130]^and_result38[131]^and_result38[132]^and_result38[133]^and_result38[134]^and_result38[135]^and_result38[136]^and_result38[137]^and_result38[138]^and_result38[139]^and_result38[140]^and_result38[141]^and_result38[142]^and_result38[143]^and_result38[144]^and_result38[145]^and_result38[146]^and_result38[147]^and_result38[148]^and_result38[149]^and_result38[150]^and_result38[151]^and_result38[152]^and_result38[153]^and_result38[154]^and_result38[155]^and_result38[156]^and_result38[157]^and_result38[158]^and_result38[159]^and_result38[160]^and_result38[161]^and_result38[162]^and_result38[163]^and_result38[164]^and_result38[165]^and_result38[166]^and_result38[167]^and_result38[168]^and_result38[169]^and_result38[170]^and_result38[171]^and_result38[172]^and_result38[173]^and_result38[174]^and_result38[175]^and_result38[176]^and_result38[177]^and_result38[178]^and_result38[179]^and_result38[180]^and_result38[181]^and_result38[182]^and_result38[183]^and_result38[184]^and_result38[185]^and_result38[186]^and_result38[187]^and_result38[188]^and_result38[189]^and_result38[190]^and_result38[191]^and_result38[192]^and_result38[193]^and_result38[194]^and_result38[195]^and_result38[196]^and_result38[197]^and_result38[198]^and_result38[199]^and_result38[200]^and_result38[201]^and_result38[202]^and_result38[203]^and_result38[204]^and_result38[205]^and_result38[206]^and_result38[207]^and_result38[208]^and_result38[209]^and_result38[210]^and_result38[211]^and_result38[212]^and_result38[213]^and_result38[214]^and_result38[215]^and_result38[216]^and_result38[217]^and_result38[218]^and_result38[219]^and_result38[220]^and_result38[221]^and_result38[222]^and_result38[223]^and_result38[224]^and_result38[225]^and_result38[226]^and_result38[227]^and_result38[228]^and_result38[229]^and_result38[230]^and_result38[231]^and_result38[232]^and_result38[233]^and_result38[234]^and_result38[235]^and_result38[236]^and_result38[237]^and_result38[238]^and_result38[239]^and_result38[240]^and_result38[241]^and_result38[242]^and_result38[243]^and_result38[244]^and_result38[245]^and_result38[246]^and_result38[247]^and_result38[248]^and_result38[249]^and_result38[250]^and_result38[251]^and_result38[252]^and_result38[253]^and_result38[254];
assign key[39]=and_result39[0]^and_result39[1]^and_result39[2]^and_result39[3]^and_result39[4]^and_result39[5]^and_result39[6]^and_result39[7]^and_result39[8]^and_result39[9]^and_result39[10]^and_result39[11]^and_result39[12]^and_result39[13]^and_result39[14]^and_result39[15]^and_result39[16]^and_result39[17]^and_result39[18]^and_result39[19]^and_result39[20]^and_result39[21]^and_result39[22]^and_result39[23]^and_result39[24]^and_result39[25]^and_result39[26]^and_result39[27]^and_result39[28]^and_result39[29]^and_result39[30]^and_result39[31]^and_result39[32]^and_result39[33]^and_result39[34]^and_result39[35]^and_result39[36]^and_result39[37]^and_result39[38]^and_result39[39]^and_result39[40]^and_result39[41]^and_result39[42]^and_result39[43]^and_result39[44]^and_result39[45]^and_result39[46]^and_result39[47]^and_result39[48]^and_result39[49]^and_result39[50]^and_result39[51]^and_result39[52]^and_result39[53]^and_result39[54]^and_result39[55]^and_result39[56]^and_result39[57]^and_result39[58]^and_result39[59]^and_result39[60]^and_result39[61]^and_result39[62]^and_result39[63]^and_result39[64]^and_result39[65]^and_result39[66]^and_result39[67]^and_result39[68]^and_result39[69]^and_result39[70]^and_result39[71]^and_result39[72]^and_result39[73]^and_result39[74]^and_result39[75]^and_result39[76]^and_result39[77]^and_result39[78]^and_result39[79]^and_result39[80]^and_result39[81]^and_result39[82]^and_result39[83]^and_result39[84]^and_result39[85]^and_result39[86]^and_result39[87]^and_result39[88]^and_result39[89]^and_result39[90]^and_result39[91]^and_result39[92]^and_result39[93]^and_result39[94]^and_result39[95]^and_result39[96]^and_result39[97]^and_result39[98]^and_result39[99]^and_result39[100]^and_result39[101]^and_result39[102]^and_result39[103]^and_result39[104]^and_result39[105]^and_result39[106]^and_result39[107]^and_result39[108]^and_result39[109]^and_result39[110]^and_result39[111]^and_result39[112]^and_result39[113]^and_result39[114]^and_result39[115]^and_result39[116]^and_result39[117]^and_result39[118]^and_result39[119]^and_result39[120]^and_result39[121]^and_result39[122]^and_result39[123]^and_result39[124]^and_result39[125]^and_result39[126]^and_result39[127]^and_result39[128]^and_result39[129]^and_result39[130]^and_result39[131]^and_result39[132]^and_result39[133]^and_result39[134]^and_result39[135]^and_result39[136]^and_result39[137]^and_result39[138]^and_result39[139]^and_result39[140]^and_result39[141]^and_result39[142]^and_result39[143]^and_result39[144]^and_result39[145]^and_result39[146]^and_result39[147]^and_result39[148]^and_result39[149]^and_result39[150]^and_result39[151]^and_result39[152]^and_result39[153]^and_result39[154]^and_result39[155]^and_result39[156]^and_result39[157]^and_result39[158]^and_result39[159]^and_result39[160]^and_result39[161]^and_result39[162]^and_result39[163]^and_result39[164]^and_result39[165]^and_result39[166]^and_result39[167]^and_result39[168]^and_result39[169]^and_result39[170]^and_result39[171]^and_result39[172]^and_result39[173]^and_result39[174]^and_result39[175]^and_result39[176]^and_result39[177]^and_result39[178]^and_result39[179]^and_result39[180]^and_result39[181]^and_result39[182]^and_result39[183]^and_result39[184]^and_result39[185]^and_result39[186]^and_result39[187]^and_result39[188]^and_result39[189]^and_result39[190]^and_result39[191]^and_result39[192]^and_result39[193]^and_result39[194]^and_result39[195]^and_result39[196]^and_result39[197]^and_result39[198]^and_result39[199]^and_result39[200]^and_result39[201]^and_result39[202]^and_result39[203]^and_result39[204]^and_result39[205]^and_result39[206]^and_result39[207]^and_result39[208]^and_result39[209]^and_result39[210]^and_result39[211]^and_result39[212]^and_result39[213]^and_result39[214]^and_result39[215]^and_result39[216]^and_result39[217]^and_result39[218]^and_result39[219]^and_result39[220]^and_result39[221]^and_result39[222]^and_result39[223]^and_result39[224]^and_result39[225]^and_result39[226]^and_result39[227]^and_result39[228]^and_result39[229]^and_result39[230]^and_result39[231]^and_result39[232]^and_result39[233]^and_result39[234]^and_result39[235]^and_result39[236]^and_result39[237]^and_result39[238]^and_result39[239]^and_result39[240]^and_result39[241]^and_result39[242]^and_result39[243]^and_result39[244]^and_result39[245]^and_result39[246]^and_result39[247]^and_result39[248]^and_result39[249]^and_result39[250]^and_result39[251]^and_result39[252]^and_result39[253]^and_result39[254];
assign key[40]=and_result40[0]^and_result40[1]^and_result40[2]^and_result40[3]^and_result40[4]^and_result40[5]^and_result40[6]^and_result40[7]^and_result40[8]^and_result40[9]^and_result40[10]^and_result40[11]^and_result40[12]^and_result40[13]^and_result40[14]^and_result40[15]^and_result40[16]^and_result40[17]^and_result40[18]^and_result40[19]^and_result40[20]^and_result40[21]^and_result40[22]^and_result40[23]^and_result40[24]^and_result40[25]^and_result40[26]^and_result40[27]^and_result40[28]^and_result40[29]^and_result40[30]^and_result40[31]^and_result40[32]^and_result40[33]^and_result40[34]^and_result40[35]^and_result40[36]^and_result40[37]^and_result40[38]^and_result40[39]^and_result40[40]^and_result40[41]^and_result40[42]^and_result40[43]^and_result40[44]^and_result40[45]^and_result40[46]^and_result40[47]^and_result40[48]^and_result40[49]^and_result40[50]^and_result40[51]^and_result40[52]^and_result40[53]^and_result40[54]^and_result40[55]^and_result40[56]^and_result40[57]^and_result40[58]^and_result40[59]^and_result40[60]^and_result40[61]^and_result40[62]^and_result40[63]^and_result40[64]^and_result40[65]^and_result40[66]^and_result40[67]^and_result40[68]^and_result40[69]^and_result40[70]^and_result40[71]^and_result40[72]^and_result40[73]^and_result40[74]^and_result40[75]^and_result40[76]^and_result40[77]^and_result40[78]^and_result40[79]^and_result40[80]^and_result40[81]^and_result40[82]^and_result40[83]^and_result40[84]^and_result40[85]^and_result40[86]^and_result40[87]^and_result40[88]^and_result40[89]^and_result40[90]^and_result40[91]^and_result40[92]^and_result40[93]^and_result40[94]^and_result40[95]^and_result40[96]^and_result40[97]^and_result40[98]^and_result40[99]^and_result40[100]^and_result40[101]^and_result40[102]^and_result40[103]^and_result40[104]^and_result40[105]^and_result40[106]^and_result40[107]^and_result40[108]^and_result40[109]^and_result40[110]^and_result40[111]^and_result40[112]^and_result40[113]^and_result40[114]^and_result40[115]^and_result40[116]^and_result40[117]^and_result40[118]^and_result40[119]^and_result40[120]^and_result40[121]^and_result40[122]^and_result40[123]^and_result40[124]^and_result40[125]^and_result40[126]^and_result40[127]^and_result40[128]^and_result40[129]^and_result40[130]^and_result40[131]^and_result40[132]^and_result40[133]^and_result40[134]^and_result40[135]^and_result40[136]^and_result40[137]^and_result40[138]^and_result40[139]^and_result40[140]^and_result40[141]^and_result40[142]^and_result40[143]^and_result40[144]^and_result40[145]^and_result40[146]^and_result40[147]^and_result40[148]^and_result40[149]^and_result40[150]^and_result40[151]^and_result40[152]^and_result40[153]^and_result40[154]^and_result40[155]^and_result40[156]^and_result40[157]^and_result40[158]^and_result40[159]^and_result40[160]^and_result40[161]^and_result40[162]^and_result40[163]^and_result40[164]^and_result40[165]^and_result40[166]^and_result40[167]^and_result40[168]^and_result40[169]^and_result40[170]^and_result40[171]^and_result40[172]^and_result40[173]^and_result40[174]^and_result40[175]^and_result40[176]^and_result40[177]^and_result40[178]^and_result40[179]^and_result40[180]^and_result40[181]^and_result40[182]^and_result40[183]^and_result40[184]^and_result40[185]^and_result40[186]^and_result40[187]^and_result40[188]^and_result40[189]^and_result40[190]^and_result40[191]^and_result40[192]^and_result40[193]^and_result40[194]^and_result40[195]^and_result40[196]^and_result40[197]^and_result40[198]^and_result40[199]^and_result40[200]^and_result40[201]^and_result40[202]^and_result40[203]^and_result40[204]^and_result40[205]^and_result40[206]^and_result40[207]^and_result40[208]^and_result40[209]^and_result40[210]^and_result40[211]^and_result40[212]^and_result40[213]^and_result40[214]^and_result40[215]^and_result40[216]^and_result40[217]^and_result40[218]^and_result40[219]^and_result40[220]^and_result40[221]^and_result40[222]^and_result40[223]^and_result40[224]^and_result40[225]^and_result40[226]^and_result40[227]^and_result40[228]^and_result40[229]^and_result40[230]^and_result40[231]^and_result40[232]^and_result40[233]^and_result40[234]^and_result40[235]^and_result40[236]^and_result40[237]^and_result40[238]^and_result40[239]^and_result40[240]^and_result40[241]^and_result40[242]^and_result40[243]^and_result40[244]^and_result40[245]^and_result40[246]^and_result40[247]^and_result40[248]^and_result40[249]^and_result40[250]^and_result40[251]^and_result40[252]^and_result40[253]^and_result40[254];
assign key[41]=and_result41[0]^and_result41[1]^and_result41[2]^and_result41[3]^and_result41[4]^and_result41[5]^and_result41[6]^and_result41[7]^and_result41[8]^and_result41[9]^and_result41[10]^and_result41[11]^and_result41[12]^and_result41[13]^and_result41[14]^and_result41[15]^and_result41[16]^and_result41[17]^and_result41[18]^and_result41[19]^and_result41[20]^and_result41[21]^and_result41[22]^and_result41[23]^and_result41[24]^and_result41[25]^and_result41[26]^and_result41[27]^and_result41[28]^and_result41[29]^and_result41[30]^and_result41[31]^and_result41[32]^and_result41[33]^and_result41[34]^and_result41[35]^and_result41[36]^and_result41[37]^and_result41[38]^and_result41[39]^and_result41[40]^and_result41[41]^and_result41[42]^and_result41[43]^and_result41[44]^and_result41[45]^and_result41[46]^and_result41[47]^and_result41[48]^and_result41[49]^and_result41[50]^and_result41[51]^and_result41[52]^and_result41[53]^and_result41[54]^and_result41[55]^and_result41[56]^and_result41[57]^and_result41[58]^and_result41[59]^and_result41[60]^and_result41[61]^and_result41[62]^and_result41[63]^and_result41[64]^and_result41[65]^and_result41[66]^and_result41[67]^and_result41[68]^and_result41[69]^and_result41[70]^and_result41[71]^and_result41[72]^and_result41[73]^and_result41[74]^and_result41[75]^and_result41[76]^and_result41[77]^and_result41[78]^and_result41[79]^and_result41[80]^and_result41[81]^and_result41[82]^and_result41[83]^and_result41[84]^and_result41[85]^and_result41[86]^and_result41[87]^and_result41[88]^and_result41[89]^and_result41[90]^and_result41[91]^and_result41[92]^and_result41[93]^and_result41[94]^and_result41[95]^and_result41[96]^and_result41[97]^and_result41[98]^and_result41[99]^and_result41[100]^and_result41[101]^and_result41[102]^and_result41[103]^and_result41[104]^and_result41[105]^and_result41[106]^and_result41[107]^and_result41[108]^and_result41[109]^and_result41[110]^and_result41[111]^and_result41[112]^and_result41[113]^and_result41[114]^and_result41[115]^and_result41[116]^and_result41[117]^and_result41[118]^and_result41[119]^and_result41[120]^and_result41[121]^and_result41[122]^and_result41[123]^and_result41[124]^and_result41[125]^and_result41[126]^and_result41[127]^and_result41[128]^and_result41[129]^and_result41[130]^and_result41[131]^and_result41[132]^and_result41[133]^and_result41[134]^and_result41[135]^and_result41[136]^and_result41[137]^and_result41[138]^and_result41[139]^and_result41[140]^and_result41[141]^and_result41[142]^and_result41[143]^and_result41[144]^and_result41[145]^and_result41[146]^and_result41[147]^and_result41[148]^and_result41[149]^and_result41[150]^and_result41[151]^and_result41[152]^and_result41[153]^and_result41[154]^and_result41[155]^and_result41[156]^and_result41[157]^and_result41[158]^and_result41[159]^and_result41[160]^and_result41[161]^and_result41[162]^and_result41[163]^and_result41[164]^and_result41[165]^and_result41[166]^and_result41[167]^and_result41[168]^and_result41[169]^and_result41[170]^and_result41[171]^and_result41[172]^and_result41[173]^and_result41[174]^and_result41[175]^and_result41[176]^and_result41[177]^and_result41[178]^and_result41[179]^and_result41[180]^and_result41[181]^and_result41[182]^and_result41[183]^and_result41[184]^and_result41[185]^and_result41[186]^and_result41[187]^and_result41[188]^and_result41[189]^and_result41[190]^and_result41[191]^and_result41[192]^and_result41[193]^and_result41[194]^and_result41[195]^and_result41[196]^and_result41[197]^and_result41[198]^and_result41[199]^and_result41[200]^and_result41[201]^and_result41[202]^and_result41[203]^and_result41[204]^and_result41[205]^and_result41[206]^and_result41[207]^and_result41[208]^and_result41[209]^and_result41[210]^and_result41[211]^and_result41[212]^and_result41[213]^and_result41[214]^and_result41[215]^and_result41[216]^and_result41[217]^and_result41[218]^and_result41[219]^and_result41[220]^and_result41[221]^and_result41[222]^and_result41[223]^and_result41[224]^and_result41[225]^and_result41[226]^and_result41[227]^and_result41[228]^and_result41[229]^and_result41[230]^and_result41[231]^and_result41[232]^and_result41[233]^and_result41[234]^and_result41[235]^and_result41[236]^and_result41[237]^and_result41[238]^and_result41[239]^and_result41[240]^and_result41[241]^and_result41[242]^and_result41[243]^and_result41[244]^and_result41[245]^and_result41[246]^and_result41[247]^and_result41[248]^and_result41[249]^and_result41[250]^and_result41[251]^and_result41[252]^and_result41[253]^and_result41[254];
assign key[42]=and_result42[0]^and_result42[1]^and_result42[2]^and_result42[3]^and_result42[4]^and_result42[5]^and_result42[6]^and_result42[7]^and_result42[8]^and_result42[9]^and_result42[10]^and_result42[11]^and_result42[12]^and_result42[13]^and_result42[14]^and_result42[15]^and_result42[16]^and_result42[17]^and_result42[18]^and_result42[19]^and_result42[20]^and_result42[21]^and_result42[22]^and_result42[23]^and_result42[24]^and_result42[25]^and_result42[26]^and_result42[27]^and_result42[28]^and_result42[29]^and_result42[30]^and_result42[31]^and_result42[32]^and_result42[33]^and_result42[34]^and_result42[35]^and_result42[36]^and_result42[37]^and_result42[38]^and_result42[39]^and_result42[40]^and_result42[41]^and_result42[42]^and_result42[43]^and_result42[44]^and_result42[45]^and_result42[46]^and_result42[47]^and_result42[48]^and_result42[49]^and_result42[50]^and_result42[51]^and_result42[52]^and_result42[53]^and_result42[54]^and_result42[55]^and_result42[56]^and_result42[57]^and_result42[58]^and_result42[59]^and_result42[60]^and_result42[61]^and_result42[62]^and_result42[63]^and_result42[64]^and_result42[65]^and_result42[66]^and_result42[67]^and_result42[68]^and_result42[69]^and_result42[70]^and_result42[71]^and_result42[72]^and_result42[73]^and_result42[74]^and_result42[75]^and_result42[76]^and_result42[77]^and_result42[78]^and_result42[79]^and_result42[80]^and_result42[81]^and_result42[82]^and_result42[83]^and_result42[84]^and_result42[85]^and_result42[86]^and_result42[87]^and_result42[88]^and_result42[89]^and_result42[90]^and_result42[91]^and_result42[92]^and_result42[93]^and_result42[94]^and_result42[95]^and_result42[96]^and_result42[97]^and_result42[98]^and_result42[99]^and_result42[100]^and_result42[101]^and_result42[102]^and_result42[103]^and_result42[104]^and_result42[105]^and_result42[106]^and_result42[107]^and_result42[108]^and_result42[109]^and_result42[110]^and_result42[111]^and_result42[112]^and_result42[113]^and_result42[114]^and_result42[115]^and_result42[116]^and_result42[117]^and_result42[118]^and_result42[119]^and_result42[120]^and_result42[121]^and_result42[122]^and_result42[123]^and_result42[124]^and_result42[125]^and_result42[126]^and_result42[127]^and_result42[128]^and_result42[129]^and_result42[130]^and_result42[131]^and_result42[132]^and_result42[133]^and_result42[134]^and_result42[135]^and_result42[136]^and_result42[137]^and_result42[138]^and_result42[139]^and_result42[140]^and_result42[141]^and_result42[142]^and_result42[143]^and_result42[144]^and_result42[145]^and_result42[146]^and_result42[147]^and_result42[148]^and_result42[149]^and_result42[150]^and_result42[151]^and_result42[152]^and_result42[153]^and_result42[154]^and_result42[155]^and_result42[156]^and_result42[157]^and_result42[158]^and_result42[159]^and_result42[160]^and_result42[161]^and_result42[162]^and_result42[163]^and_result42[164]^and_result42[165]^and_result42[166]^and_result42[167]^and_result42[168]^and_result42[169]^and_result42[170]^and_result42[171]^and_result42[172]^and_result42[173]^and_result42[174]^and_result42[175]^and_result42[176]^and_result42[177]^and_result42[178]^and_result42[179]^and_result42[180]^and_result42[181]^and_result42[182]^and_result42[183]^and_result42[184]^and_result42[185]^and_result42[186]^and_result42[187]^and_result42[188]^and_result42[189]^and_result42[190]^and_result42[191]^and_result42[192]^and_result42[193]^and_result42[194]^and_result42[195]^and_result42[196]^and_result42[197]^and_result42[198]^and_result42[199]^and_result42[200]^and_result42[201]^and_result42[202]^and_result42[203]^and_result42[204]^and_result42[205]^and_result42[206]^and_result42[207]^and_result42[208]^and_result42[209]^and_result42[210]^and_result42[211]^and_result42[212]^and_result42[213]^and_result42[214]^and_result42[215]^and_result42[216]^and_result42[217]^and_result42[218]^and_result42[219]^and_result42[220]^and_result42[221]^and_result42[222]^and_result42[223]^and_result42[224]^and_result42[225]^and_result42[226]^and_result42[227]^and_result42[228]^and_result42[229]^and_result42[230]^and_result42[231]^and_result42[232]^and_result42[233]^and_result42[234]^and_result42[235]^and_result42[236]^and_result42[237]^and_result42[238]^and_result42[239]^and_result42[240]^and_result42[241]^and_result42[242]^and_result42[243]^and_result42[244]^and_result42[245]^and_result42[246]^and_result42[247]^and_result42[248]^and_result42[249]^and_result42[250]^and_result42[251]^and_result42[252]^and_result42[253]^and_result42[254];
assign key[43]=and_result43[0]^and_result43[1]^and_result43[2]^and_result43[3]^and_result43[4]^and_result43[5]^and_result43[6]^and_result43[7]^and_result43[8]^and_result43[9]^and_result43[10]^and_result43[11]^and_result43[12]^and_result43[13]^and_result43[14]^and_result43[15]^and_result43[16]^and_result43[17]^and_result43[18]^and_result43[19]^and_result43[20]^and_result43[21]^and_result43[22]^and_result43[23]^and_result43[24]^and_result43[25]^and_result43[26]^and_result43[27]^and_result43[28]^and_result43[29]^and_result43[30]^and_result43[31]^and_result43[32]^and_result43[33]^and_result43[34]^and_result43[35]^and_result43[36]^and_result43[37]^and_result43[38]^and_result43[39]^and_result43[40]^and_result43[41]^and_result43[42]^and_result43[43]^and_result43[44]^and_result43[45]^and_result43[46]^and_result43[47]^and_result43[48]^and_result43[49]^and_result43[50]^and_result43[51]^and_result43[52]^and_result43[53]^and_result43[54]^and_result43[55]^and_result43[56]^and_result43[57]^and_result43[58]^and_result43[59]^and_result43[60]^and_result43[61]^and_result43[62]^and_result43[63]^and_result43[64]^and_result43[65]^and_result43[66]^and_result43[67]^and_result43[68]^and_result43[69]^and_result43[70]^and_result43[71]^and_result43[72]^and_result43[73]^and_result43[74]^and_result43[75]^and_result43[76]^and_result43[77]^and_result43[78]^and_result43[79]^and_result43[80]^and_result43[81]^and_result43[82]^and_result43[83]^and_result43[84]^and_result43[85]^and_result43[86]^and_result43[87]^and_result43[88]^and_result43[89]^and_result43[90]^and_result43[91]^and_result43[92]^and_result43[93]^and_result43[94]^and_result43[95]^and_result43[96]^and_result43[97]^and_result43[98]^and_result43[99]^and_result43[100]^and_result43[101]^and_result43[102]^and_result43[103]^and_result43[104]^and_result43[105]^and_result43[106]^and_result43[107]^and_result43[108]^and_result43[109]^and_result43[110]^and_result43[111]^and_result43[112]^and_result43[113]^and_result43[114]^and_result43[115]^and_result43[116]^and_result43[117]^and_result43[118]^and_result43[119]^and_result43[120]^and_result43[121]^and_result43[122]^and_result43[123]^and_result43[124]^and_result43[125]^and_result43[126]^and_result43[127]^and_result43[128]^and_result43[129]^and_result43[130]^and_result43[131]^and_result43[132]^and_result43[133]^and_result43[134]^and_result43[135]^and_result43[136]^and_result43[137]^and_result43[138]^and_result43[139]^and_result43[140]^and_result43[141]^and_result43[142]^and_result43[143]^and_result43[144]^and_result43[145]^and_result43[146]^and_result43[147]^and_result43[148]^and_result43[149]^and_result43[150]^and_result43[151]^and_result43[152]^and_result43[153]^and_result43[154]^and_result43[155]^and_result43[156]^and_result43[157]^and_result43[158]^and_result43[159]^and_result43[160]^and_result43[161]^and_result43[162]^and_result43[163]^and_result43[164]^and_result43[165]^and_result43[166]^and_result43[167]^and_result43[168]^and_result43[169]^and_result43[170]^and_result43[171]^and_result43[172]^and_result43[173]^and_result43[174]^and_result43[175]^and_result43[176]^and_result43[177]^and_result43[178]^and_result43[179]^and_result43[180]^and_result43[181]^and_result43[182]^and_result43[183]^and_result43[184]^and_result43[185]^and_result43[186]^and_result43[187]^and_result43[188]^and_result43[189]^and_result43[190]^and_result43[191]^and_result43[192]^and_result43[193]^and_result43[194]^and_result43[195]^and_result43[196]^and_result43[197]^and_result43[198]^and_result43[199]^and_result43[200]^and_result43[201]^and_result43[202]^and_result43[203]^and_result43[204]^and_result43[205]^and_result43[206]^and_result43[207]^and_result43[208]^and_result43[209]^and_result43[210]^and_result43[211]^and_result43[212]^and_result43[213]^and_result43[214]^and_result43[215]^and_result43[216]^and_result43[217]^and_result43[218]^and_result43[219]^and_result43[220]^and_result43[221]^and_result43[222]^and_result43[223]^and_result43[224]^and_result43[225]^and_result43[226]^and_result43[227]^and_result43[228]^and_result43[229]^and_result43[230]^and_result43[231]^and_result43[232]^and_result43[233]^and_result43[234]^and_result43[235]^and_result43[236]^and_result43[237]^and_result43[238]^and_result43[239]^and_result43[240]^and_result43[241]^and_result43[242]^and_result43[243]^and_result43[244]^and_result43[245]^and_result43[246]^and_result43[247]^and_result43[248]^and_result43[249]^and_result43[250]^and_result43[251]^and_result43[252]^and_result43[253]^and_result43[254];
assign key[44]=and_result44[0]^and_result44[1]^and_result44[2]^and_result44[3]^and_result44[4]^and_result44[5]^and_result44[6]^and_result44[7]^and_result44[8]^and_result44[9]^and_result44[10]^and_result44[11]^and_result44[12]^and_result44[13]^and_result44[14]^and_result44[15]^and_result44[16]^and_result44[17]^and_result44[18]^and_result44[19]^and_result44[20]^and_result44[21]^and_result44[22]^and_result44[23]^and_result44[24]^and_result44[25]^and_result44[26]^and_result44[27]^and_result44[28]^and_result44[29]^and_result44[30]^and_result44[31]^and_result44[32]^and_result44[33]^and_result44[34]^and_result44[35]^and_result44[36]^and_result44[37]^and_result44[38]^and_result44[39]^and_result44[40]^and_result44[41]^and_result44[42]^and_result44[43]^and_result44[44]^and_result44[45]^and_result44[46]^and_result44[47]^and_result44[48]^and_result44[49]^and_result44[50]^and_result44[51]^and_result44[52]^and_result44[53]^and_result44[54]^and_result44[55]^and_result44[56]^and_result44[57]^and_result44[58]^and_result44[59]^and_result44[60]^and_result44[61]^and_result44[62]^and_result44[63]^and_result44[64]^and_result44[65]^and_result44[66]^and_result44[67]^and_result44[68]^and_result44[69]^and_result44[70]^and_result44[71]^and_result44[72]^and_result44[73]^and_result44[74]^and_result44[75]^and_result44[76]^and_result44[77]^and_result44[78]^and_result44[79]^and_result44[80]^and_result44[81]^and_result44[82]^and_result44[83]^and_result44[84]^and_result44[85]^and_result44[86]^and_result44[87]^and_result44[88]^and_result44[89]^and_result44[90]^and_result44[91]^and_result44[92]^and_result44[93]^and_result44[94]^and_result44[95]^and_result44[96]^and_result44[97]^and_result44[98]^and_result44[99]^and_result44[100]^and_result44[101]^and_result44[102]^and_result44[103]^and_result44[104]^and_result44[105]^and_result44[106]^and_result44[107]^and_result44[108]^and_result44[109]^and_result44[110]^and_result44[111]^and_result44[112]^and_result44[113]^and_result44[114]^and_result44[115]^and_result44[116]^and_result44[117]^and_result44[118]^and_result44[119]^and_result44[120]^and_result44[121]^and_result44[122]^and_result44[123]^and_result44[124]^and_result44[125]^and_result44[126]^and_result44[127]^and_result44[128]^and_result44[129]^and_result44[130]^and_result44[131]^and_result44[132]^and_result44[133]^and_result44[134]^and_result44[135]^and_result44[136]^and_result44[137]^and_result44[138]^and_result44[139]^and_result44[140]^and_result44[141]^and_result44[142]^and_result44[143]^and_result44[144]^and_result44[145]^and_result44[146]^and_result44[147]^and_result44[148]^and_result44[149]^and_result44[150]^and_result44[151]^and_result44[152]^and_result44[153]^and_result44[154]^and_result44[155]^and_result44[156]^and_result44[157]^and_result44[158]^and_result44[159]^and_result44[160]^and_result44[161]^and_result44[162]^and_result44[163]^and_result44[164]^and_result44[165]^and_result44[166]^and_result44[167]^and_result44[168]^and_result44[169]^and_result44[170]^and_result44[171]^and_result44[172]^and_result44[173]^and_result44[174]^and_result44[175]^and_result44[176]^and_result44[177]^and_result44[178]^and_result44[179]^and_result44[180]^and_result44[181]^and_result44[182]^and_result44[183]^and_result44[184]^and_result44[185]^and_result44[186]^and_result44[187]^and_result44[188]^and_result44[189]^and_result44[190]^and_result44[191]^and_result44[192]^and_result44[193]^and_result44[194]^and_result44[195]^and_result44[196]^and_result44[197]^and_result44[198]^and_result44[199]^and_result44[200]^and_result44[201]^and_result44[202]^and_result44[203]^and_result44[204]^and_result44[205]^and_result44[206]^and_result44[207]^and_result44[208]^and_result44[209]^and_result44[210]^and_result44[211]^and_result44[212]^and_result44[213]^and_result44[214]^and_result44[215]^and_result44[216]^and_result44[217]^and_result44[218]^and_result44[219]^and_result44[220]^and_result44[221]^and_result44[222]^and_result44[223]^and_result44[224]^and_result44[225]^and_result44[226]^and_result44[227]^and_result44[228]^and_result44[229]^and_result44[230]^and_result44[231]^and_result44[232]^and_result44[233]^and_result44[234]^and_result44[235]^and_result44[236]^and_result44[237]^and_result44[238]^and_result44[239]^and_result44[240]^and_result44[241]^and_result44[242]^and_result44[243]^and_result44[244]^and_result44[245]^and_result44[246]^and_result44[247]^and_result44[248]^and_result44[249]^and_result44[250]^and_result44[251]^and_result44[252]^and_result44[253]^and_result44[254];
assign key[45]=and_result45[0]^and_result45[1]^and_result45[2]^and_result45[3]^and_result45[4]^and_result45[5]^and_result45[6]^and_result45[7]^and_result45[8]^and_result45[9]^and_result45[10]^and_result45[11]^and_result45[12]^and_result45[13]^and_result45[14]^and_result45[15]^and_result45[16]^and_result45[17]^and_result45[18]^and_result45[19]^and_result45[20]^and_result45[21]^and_result45[22]^and_result45[23]^and_result45[24]^and_result45[25]^and_result45[26]^and_result45[27]^and_result45[28]^and_result45[29]^and_result45[30]^and_result45[31]^and_result45[32]^and_result45[33]^and_result45[34]^and_result45[35]^and_result45[36]^and_result45[37]^and_result45[38]^and_result45[39]^and_result45[40]^and_result45[41]^and_result45[42]^and_result45[43]^and_result45[44]^and_result45[45]^and_result45[46]^and_result45[47]^and_result45[48]^and_result45[49]^and_result45[50]^and_result45[51]^and_result45[52]^and_result45[53]^and_result45[54]^and_result45[55]^and_result45[56]^and_result45[57]^and_result45[58]^and_result45[59]^and_result45[60]^and_result45[61]^and_result45[62]^and_result45[63]^and_result45[64]^and_result45[65]^and_result45[66]^and_result45[67]^and_result45[68]^and_result45[69]^and_result45[70]^and_result45[71]^and_result45[72]^and_result45[73]^and_result45[74]^and_result45[75]^and_result45[76]^and_result45[77]^and_result45[78]^and_result45[79]^and_result45[80]^and_result45[81]^and_result45[82]^and_result45[83]^and_result45[84]^and_result45[85]^and_result45[86]^and_result45[87]^and_result45[88]^and_result45[89]^and_result45[90]^and_result45[91]^and_result45[92]^and_result45[93]^and_result45[94]^and_result45[95]^and_result45[96]^and_result45[97]^and_result45[98]^and_result45[99]^and_result45[100]^and_result45[101]^and_result45[102]^and_result45[103]^and_result45[104]^and_result45[105]^and_result45[106]^and_result45[107]^and_result45[108]^and_result45[109]^and_result45[110]^and_result45[111]^and_result45[112]^and_result45[113]^and_result45[114]^and_result45[115]^and_result45[116]^and_result45[117]^and_result45[118]^and_result45[119]^and_result45[120]^and_result45[121]^and_result45[122]^and_result45[123]^and_result45[124]^and_result45[125]^and_result45[126]^and_result45[127]^and_result45[128]^and_result45[129]^and_result45[130]^and_result45[131]^and_result45[132]^and_result45[133]^and_result45[134]^and_result45[135]^and_result45[136]^and_result45[137]^and_result45[138]^and_result45[139]^and_result45[140]^and_result45[141]^and_result45[142]^and_result45[143]^and_result45[144]^and_result45[145]^and_result45[146]^and_result45[147]^and_result45[148]^and_result45[149]^and_result45[150]^and_result45[151]^and_result45[152]^and_result45[153]^and_result45[154]^and_result45[155]^and_result45[156]^and_result45[157]^and_result45[158]^and_result45[159]^and_result45[160]^and_result45[161]^and_result45[162]^and_result45[163]^and_result45[164]^and_result45[165]^and_result45[166]^and_result45[167]^and_result45[168]^and_result45[169]^and_result45[170]^and_result45[171]^and_result45[172]^and_result45[173]^and_result45[174]^and_result45[175]^and_result45[176]^and_result45[177]^and_result45[178]^and_result45[179]^and_result45[180]^and_result45[181]^and_result45[182]^and_result45[183]^and_result45[184]^and_result45[185]^and_result45[186]^and_result45[187]^and_result45[188]^and_result45[189]^and_result45[190]^and_result45[191]^and_result45[192]^and_result45[193]^and_result45[194]^and_result45[195]^and_result45[196]^and_result45[197]^and_result45[198]^and_result45[199]^and_result45[200]^and_result45[201]^and_result45[202]^and_result45[203]^and_result45[204]^and_result45[205]^and_result45[206]^and_result45[207]^and_result45[208]^and_result45[209]^and_result45[210]^and_result45[211]^and_result45[212]^and_result45[213]^and_result45[214]^and_result45[215]^and_result45[216]^and_result45[217]^and_result45[218]^and_result45[219]^and_result45[220]^and_result45[221]^and_result45[222]^and_result45[223]^and_result45[224]^and_result45[225]^and_result45[226]^and_result45[227]^and_result45[228]^and_result45[229]^and_result45[230]^and_result45[231]^and_result45[232]^and_result45[233]^and_result45[234]^and_result45[235]^and_result45[236]^and_result45[237]^and_result45[238]^and_result45[239]^and_result45[240]^and_result45[241]^and_result45[242]^and_result45[243]^and_result45[244]^and_result45[245]^and_result45[246]^and_result45[247]^and_result45[248]^and_result45[249]^and_result45[250]^and_result45[251]^and_result45[252]^and_result45[253]^and_result45[254];
assign key[46]=and_result46[0]^and_result46[1]^and_result46[2]^and_result46[3]^and_result46[4]^and_result46[5]^and_result46[6]^and_result46[7]^and_result46[8]^and_result46[9]^and_result46[10]^and_result46[11]^and_result46[12]^and_result46[13]^and_result46[14]^and_result46[15]^and_result46[16]^and_result46[17]^and_result46[18]^and_result46[19]^and_result46[20]^and_result46[21]^and_result46[22]^and_result46[23]^and_result46[24]^and_result46[25]^and_result46[26]^and_result46[27]^and_result46[28]^and_result46[29]^and_result46[30]^and_result46[31]^and_result46[32]^and_result46[33]^and_result46[34]^and_result46[35]^and_result46[36]^and_result46[37]^and_result46[38]^and_result46[39]^and_result46[40]^and_result46[41]^and_result46[42]^and_result46[43]^and_result46[44]^and_result46[45]^and_result46[46]^and_result46[47]^and_result46[48]^and_result46[49]^and_result46[50]^and_result46[51]^and_result46[52]^and_result46[53]^and_result46[54]^and_result46[55]^and_result46[56]^and_result46[57]^and_result46[58]^and_result46[59]^and_result46[60]^and_result46[61]^and_result46[62]^and_result46[63]^and_result46[64]^and_result46[65]^and_result46[66]^and_result46[67]^and_result46[68]^and_result46[69]^and_result46[70]^and_result46[71]^and_result46[72]^and_result46[73]^and_result46[74]^and_result46[75]^and_result46[76]^and_result46[77]^and_result46[78]^and_result46[79]^and_result46[80]^and_result46[81]^and_result46[82]^and_result46[83]^and_result46[84]^and_result46[85]^and_result46[86]^and_result46[87]^and_result46[88]^and_result46[89]^and_result46[90]^and_result46[91]^and_result46[92]^and_result46[93]^and_result46[94]^and_result46[95]^and_result46[96]^and_result46[97]^and_result46[98]^and_result46[99]^and_result46[100]^and_result46[101]^and_result46[102]^and_result46[103]^and_result46[104]^and_result46[105]^and_result46[106]^and_result46[107]^and_result46[108]^and_result46[109]^and_result46[110]^and_result46[111]^and_result46[112]^and_result46[113]^and_result46[114]^and_result46[115]^and_result46[116]^and_result46[117]^and_result46[118]^and_result46[119]^and_result46[120]^and_result46[121]^and_result46[122]^and_result46[123]^and_result46[124]^and_result46[125]^and_result46[126]^and_result46[127]^and_result46[128]^and_result46[129]^and_result46[130]^and_result46[131]^and_result46[132]^and_result46[133]^and_result46[134]^and_result46[135]^and_result46[136]^and_result46[137]^and_result46[138]^and_result46[139]^and_result46[140]^and_result46[141]^and_result46[142]^and_result46[143]^and_result46[144]^and_result46[145]^and_result46[146]^and_result46[147]^and_result46[148]^and_result46[149]^and_result46[150]^and_result46[151]^and_result46[152]^and_result46[153]^and_result46[154]^and_result46[155]^and_result46[156]^and_result46[157]^and_result46[158]^and_result46[159]^and_result46[160]^and_result46[161]^and_result46[162]^and_result46[163]^and_result46[164]^and_result46[165]^and_result46[166]^and_result46[167]^and_result46[168]^and_result46[169]^and_result46[170]^and_result46[171]^and_result46[172]^and_result46[173]^and_result46[174]^and_result46[175]^and_result46[176]^and_result46[177]^and_result46[178]^and_result46[179]^and_result46[180]^and_result46[181]^and_result46[182]^and_result46[183]^and_result46[184]^and_result46[185]^and_result46[186]^and_result46[187]^and_result46[188]^and_result46[189]^and_result46[190]^and_result46[191]^and_result46[192]^and_result46[193]^and_result46[194]^and_result46[195]^and_result46[196]^and_result46[197]^and_result46[198]^and_result46[199]^and_result46[200]^and_result46[201]^and_result46[202]^and_result46[203]^and_result46[204]^and_result46[205]^and_result46[206]^and_result46[207]^and_result46[208]^and_result46[209]^and_result46[210]^and_result46[211]^and_result46[212]^and_result46[213]^and_result46[214]^and_result46[215]^and_result46[216]^and_result46[217]^and_result46[218]^and_result46[219]^and_result46[220]^and_result46[221]^and_result46[222]^and_result46[223]^and_result46[224]^and_result46[225]^and_result46[226]^and_result46[227]^and_result46[228]^and_result46[229]^and_result46[230]^and_result46[231]^and_result46[232]^and_result46[233]^and_result46[234]^and_result46[235]^and_result46[236]^and_result46[237]^and_result46[238]^and_result46[239]^and_result46[240]^and_result46[241]^and_result46[242]^and_result46[243]^and_result46[244]^and_result46[245]^and_result46[246]^and_result46[247]^and_result46[248]^and_result46[249]^and_result46[250]^and_result46[251]^and_result46[252]^and_result46[253]^and_result46[254];
assign key[47]=and_result47[0]^and_result47[1]^and_result47[2]^and_result47[3]^and_result47[4]^and_result47[5]^and_result47[6]^and_result47[7]^and_result47[8]^and_result47[9]^and_result47[10]^and_result47[11]^and_result47[12]^and_result47[13]^and_result47[14]^and_result47[15]^and_result47[16]^and_result47[17]^and_result47[18]^and_result47[19]^and_result47[20]^and_result47[21]^and_result47[22]^and_result47[23]^and_result47[24]^and_result47[25]^and_result47[26]^and_result47[27]^and_result47[28]^and_result47[29]^and_result47[30]^and_result47[31]^and_result47[32]^and_result47[33]^and_result47[34]^and_result47[35]^and_result47[36]^and_result47[37]^and_result47[38]^and_result47[39]^and_result47[40]^and_result47[41]^and_result47[42]^and_result47[43]^and_result47[44]^and_result47[45]^and_result47[46]^and_result47[47]^and_result47[48]^and_result47[49]^and_result47[50]^and_result47[51]^and_result47[52]^and_result47[53]^and_result47[54]^and_result47[55]^and_result47[56]^and_result47[57]^and_result47[58]^and_result47[59]^and_result47[60]^and_result47[61]^and_result47[62]^and_result47[63]^and_result47[64]^and_result47[65]^and_result47[66]^and_result47[67]^and_result47[68]^and_result47[69]^and_result47[70]^and_result47[71]^and_result47[72]^and_result47[73]^and_result47[74]^and_result47[75]^and_result47[76]^and_result47[77]^and_result47[78]^and_result47[79]^and_result47[80]^and_result47[81]^and_result47[82]^and_result47[83]^and_result47[84]^and_result47[85]^and_result47[86]^and_result47[87]^and_result47[88]^and_result47[89]^and_result47[90]^and_result47[91]^and_result47[92]^and_result47[93]^and_result47[94]^and_result47[95]^and_result47[96]^and_result47[97]^and_result47[98]^and_result47[99]^and_result47[100]^and_result47[101]^and_result47[102]^and_result47[103]^and_result47[104]^and_result47[105]^and_result47[106]^and_result47[107]^and_result47[108]^and_result47[109]^and_result47[110]^and_result47[111]^and_result47[112]^and_result47[113]^and_result47[114]^and_result47[115]^and_result47[116]^and_result47[117]^and_result47[118]^and_result47[119]^and_result47[120]^and_result47[121]^and_result47[122]^and_result47[123]^and_result47[124]^and_result47[125]^and_result47[126]^and_result47[127]^and_result47[128]^and_result47[129]^and_result47[130]^and_result47[131]^and_result47[132]^and_result47[133]^and_result47[134]^and_result47[135]^and_result47[136]^and_result47[137]^and_result47[138]^and_result47[139]^and_result47[140]^and_result47[141]^and_result47[142]^and_result47[143]^and_result47[144]^and_result47[145]^and_result47[146]^and_result47[147]^and_result47[148]^and_result47[149]^and_result47[150]^and_result47[151]^and_result47[152]^and_result47[153]^and_result47[154]^and_result47[155]^and_result47[156]^and_result47[157]^and_result47[158]^and_result47[159]^and_result47[160]^and_result47[161]^and_result47[162]^and_result47[163]^and_result47[164]^and_result47[165]^and_result47[166]^and_result47[167]^and_result47[168]^and_result47[169]^and_result47[170]^and_result47[171]^and_result47[172]^and_result47[173]^and_result47[174]^and_result47[175]^and_result47[176]^and_result47[177]^and_result47[178]^and_result47[179]^and_result47[180]^and_result47[181]^and_result47[182]^and_result47[183]^and_result47[184]^and_result47[185]^and_result47[186]^and_result47[187]^and_result47[188]^and_result47[189]^and_result47[190]^and_result47[191]^and_result47[192]^and_result47[193]^and_result47[194]^and_result47[195]^and_result47[196]^and_result47[197]^and_result47[198]^and_result47[199]^and_result47[200]^and_result47[201]^and_result47[202]^and_result47[203]^and_result47[204]^and_result47[205]^and_result47[206]^and_result47[207]^and_result47[208]^and_result47[209]^and_result47[210]^and_result47[211]^and_result47[212]^and_result47[213]^and_result47[214]^and_result47[215]^and_result47[216]^and_result47[217]^and_result47[218]^and_result47[219]^and_result47[220]^and_result47[221]^and_result47[222]^and_result47[223]^and_result47[224]^and_result47[225]^and_result47[226]^and_result47[227]^and_result47[228]^and_result47[229]^and_result47[230]^and_result47[231]^and_result47[232]^and_result47[233]^and_result47[234]^and_result47[235]^and_result47[236]^and_result47[237]^and_result47[238]^and_result47[239]^and_result47[240]^and_result47[241]^and_result47[242]^and_result47[243]^and_result47[244]^and_result47[245]^and_result47[246]^and_result47[247]^and_result47[248]^and_result47[249]^and_result47[250]^and_result47[251]^and_result47[252]^and_result47[253]^and_result47[254];
assign key[48]=and_result48[0]^and_result48[1]^and_result48[2]^and_result48[3]^and_result48[4]^and_result48[5]^and_result48[6]^and_result48[7]^and_result48[8]^and_result48[9]^and_result48[10]^and_result48[11]^and_result48[12]^and_result48[13]^and_result48[14]^and_result48[15]^and_result48[16]^and_result48[17]^and_result48[18]^and_result48[19]^and_result48[20]^and_result48[21]^and_result48[22]^and_result48[23]^and_result48[24]^and_result48[25]^and_result48[26]^and_result48[27]^and_result48[28]^and_result48[29]^and_result48[30]^and_result48[31]^and_result48[32]^and_result48[33]^and_result48[34]^and_result48[35]^and_result48[36]^and_result48[37]^and_result48[38]^and_result48[39]^and_result48[40]^and_result48[41]^and_result48[42]^and_result48[43]^and_result48[44]^and_result48[45]^and_result48[46]^and_result48[47]^and_result48[48]^and_result48[49]^and_result48[50]^and_result48[51]^and_result48[52]^and_result48[53]^and_result48[54]^and_result48[55]^and_result48[56]^and_result48[57]^and_result48[58]^and_result48[59]^and_result48[60]^and_result48[61]^and_result48[62]^and_result48[63]^and_result48[64]^and_result48[65]^and_result48[66]^and_result48[67]^and_result48[68]^and_result48[69]^and_result48[70]^and_result48[71]^and_result48[72]^and_result48[73]^and_result48[74]^and_result48[75]^and_result48[76]^and_result48[77]^and_result48[78]^and_result48[79]^and_result48[80]^and_result48[81]^and_result48[82]^and_result48[83]^and_result48[84]^and_result48[85]^and_result48[86]^and_result48[87]^and_result48[88]^and_result48[89]^and_result48[90]^and_result48[91]^and_result48[92]^and_result48[93]^and_result48[94]^and_result48[95]^and_result48[96]^and_result48[97]^and_result48[98]^and_result48[99]^and_result48[100]^and_result48[101]^and_result48[102]^and_result48[103]^and_result48[104]^and_result48[105]^and_result48[106]^and_result48[107]^and_result48[108]^and_result48[109]^and_result48[110]^and_result48[111]^and_result48[112]^and_result48[113]^and_result48[114]^and_result48[115]^and_result48[116]^and_result48[117]^and_result48[118]^and_result48[119]^and_result48[120]^and_result48[121]^and_result48[122]^and_result48[123]^and_result48[124]^and_result48[125]^and_result48[126]^and_result48[127]^and_result48[128]^and_result48[129]^and_result48[130]^and_result48[131]^and_result48[132]^and_result48[133]^and_result48[134]^and_result48[135]^and_result48[136]^and_result48[137]^and_result48[138]^and_result48[139]^and_result48[140]^and_result48[141]^and_result48[142]^and_result48[143]^and_result48[144]^and_result48[145]^and_result48[146]^and_result48[147]^and_result48[148]^and_result48[149]^and_result48[150]^and_result48[151]^and_result48[152]^and_result48[153]^and_result48[154]^and_result48[155]^and_result48[156]^and_result48[157]^and_result48[158]^and_result48[159]^and_result48[160]^and_result48[161]^and_result48[162]^and_result48[163]^and_result48[164]^and_result48[165]^and_result48[166]^and_result48[167]^and_result48[168]^and_result48[169]^and_result48[170]^and_result48[171]^and_result48[172]^and_result48[173]^and_result48[174]^and_result48[175]^and_result48[176]^and_result48[177]^and_result48[178]^and_result48[179]^and_result48[180]^and_result48[181]^and_result48[182]^and_result48[183]^and_result48[184]^and_result48[185]^and_result48[186]^and_result48[187]^and_result48[188]^and_result48[189]^and_result48[190]^and_result48[191]^and_result48[192]^and_result48[193]^and_result48[194]^and_result48[195]^and_result48[196]^and_result48[197]^and_result48[198]^and_result48[199]^and_result48[200]^and_result48[201]^and_result48[202]^and_result48[203]^and_result48[204]^and_result48[205]^and_result48[206]^and_result48[207]^and_result48[208]^and_result48[209]^and_result48[210]^and_result48[211]^and_result48[212]^and_result48[213]^and_result48[214]^and_result48[215]^and_result48[216]^and_result48[217]^and_result48[218]^and_result48[219]^and_result48[220]^and_result48[221]^and_result48[222]^and_result48[223]^and_result48[224]^and_result48[225]^and_result48[226]^and_result48[227]^and_result48[228]^and_result48[229]^and_result48[230]^and_result48[231]^and_result48[232]^and_result48[233]^and_result48[234]^and_result48[235]^and_result48[236]^and_result48[237]^and_result48[238]^and_result48[239]^and_result48[240]^and_result48[241]^and_result48[242]^and_result48[243]^and_result48[244]^and_result48[245]^and_result48[246]^and_result48[247]^and_result48[248]^and_result48[249]^and_result48[250]^and_result48[251]^and_result48[252]^and_result48[253]^and_result48[254];
assign key[49]=and_result49[0]^and_result49[1]^and_result49[2]^and_result49[3]^and_result49[4]^and_result49[5]^and_result49[6]^and_result49[7]^and_result49[8]^and_result49[9]^and_result49[10]^and_result49[11]^and_result49[12]^and_result49[13]^and_result49[14]^and_result49[15]^and_result49[16]^and_result49[17]^and_result49[18]^and_result49[19]^and_result49[20]^and_result49[21]^and_result49[22]^and_result49[23]^and_result49[24]^and_result49[25]^and_result49[26]^and_result49[27]^and_result49[28]^and_result49[29]^and_result49[30]^and_result49[31]^and_result49[32]^and_result49[33]^and_result49[34]^and_result49[35]^and_result49[36]^and_result49[37]^and_result49[38]^and_result49[39]^and_result49[40]^and_result49[41]^and_result49[42]^and_result49[43]^and_result49[44]^and_result49[45]^and_result49[46]^and_result49[47]^and_result49[48]^and_result49[49]^and_result49[50]^and_result49[51]^and_result49[52]^and_result49[53]^and_result49[54]^and_result49[55]^and_result49[56]^and_result49[57]^and_result49[58]^and_result49[59]^and_result49[60]^and_result49[61]^and_result49[62]^and_result49[63]^and_result49[64]^and_result49[65]^and_result49[66]^and_result49[67]^and_result49[68]^and_result49[69]^and_result49[70]^and_result49[71]^and_result49[72]^and_result49[73]^and_result49[74]^and_result49[75]^and_result49[76]^and_result49[77]^and_result49[78]^and_result49[79]^and_result49[80]^and_result49[81]^and_result49[82]^and_result49[83]^and_result49[84]^and_result49[85]^and_result49[86]^and_result49[87]^and_result49[88]^and_result49[89]^and_result49[90]^and_result49[91]^and_result49[92]^and_result49[93]^and_result49[94]^and_result49[95]^and_result49[96]^and_result49[97]^and_result49[98]^and_result49[99]^and_result49[100]^and_result49[101]^and_result49[102]^and_result49[103]^and_result49[104]^and_result49[105]^and_result49[106]^and_result49[107]^and_result49[108]^and_result49[109]^and_result49[110]^and_result49[111]^and_result49[112]^and_result49[113]^and_result49[114]^and_result49[115]^and_result49[116]^and_result49[117]^and_result49[118]^and_result49[119]^and_result49[120]^and_result49[121]^and_result49[122]^and_result49[123]^and_result49[124]^and_result49[125]^and_result49[126]^and_result49[127]^and_result49[128]^and_result49[129]^and_result49[130]^and_result49[131]^and_result49[132]^and_result49[133]^and_result49[134]^and_result49[135]^and_result49[136]^and_result49[137]^and_result49[138]^and_result49[139]^and_result49[140]^and_result49[141]^and_result49[142]^and_result49[143]^and_result49[144]^and_result49[145]^and_result49[146]^and_result49[147]^and_result49[148]^and_result49[149]^and_result49[150]^and_result49[151]^and_result49[152]^and_result49[153]^and_result49[154]^and_result49[155]^and_result49[156]^and_result49[157]^and_result49[158]^and_result49[159]^and_result49[160]^and_result49[161]^and_result49[162]^and_result49[163]^and_result49[164]^and_result49[165]^and_result49[166]^and_result49[167]^and_result49[168]^and_result49[169]^and_result49[170]^and_result49[171]^and_result49[172]^and_result49[173]^and_result49[174]^and_result49[175]^and_result49[176]^and_result49[177]^and_result49[178]^and_result49[179]^and_result49[180]^and_result49[181]^and_result49[182]^and_result49[183]^and_result49[184]^and_result49[185]^and_result49[186]^and_result49[187]^and_result49[188]^and_result49[189]^and_result49[190]^and_result49[191]^and_result49[192]^and_result49[193]^and_result49[194]^and_result49[195]^and_result49[196]^and_result49[197]^and_result49[198]^and_result49[199]^and_result49[200]^and_result49[201]^and_result49[202]^and_result49[203]^and_result49[204]^and_result49[205]^and_result49[206]^and_result49[207]^and_result49[208]^and_result49[209]^and_result49[210]^and_result49[211]^and_result49[212]^and_result49[213]^and_result49[214]^and_result49[215]^and_result49[216]^and_result49[217]^and_result49[218]^and_result49[219]^and_result49[220]^and_result49[221]^and_result49[222]^and_result49[223]^and_result49[224]^and_result49[225]^and_result49[226]^and_result49[227]^and_result49[228]^and_result49[229]^and_result49[230]^and_result49[231]^and_result49[232]^and_result49[233]^and_result49[234]^and_result49[235]^and_result49[236]^and_result49[237]^and_result49[238]^and_result49[239]^and_result49[240]^and_result49[241]^and_result49[242]^and_result49[243]^and_result49[244]^and_result49[245]^and_result49[246]^and_result49[247]^and_result49[248]^and_result49[249]^and_result49[250]^and_result49[251]^and_result49[252]^and_result49[253]^and_result49[254];
assign key[50]=and_result50[0]^and_result50[1]^and_result50[2]^and_result50[3]^and_result50[4]^and_result50[5]^and_result50[6]^and_result50[7]^and_result50[8]^and_result50[9]^and_result50[10]^and_result50[11]^and_result50[12]^and_result50[13]^and_result50[14]^and_result50[15]^and_result50[16]^and_result50[17]^and_result50[18]^and_result50[19]^and_result50[20]^and_result50[21]^and_result50[22]^and_result50[23]^and_result50[24]^and_result50[25]^and_result50[26]^and_result50[27]^and_result50[28]^and_result50[29]^and_result50[30]^and_result50[31]^and_result50[32]^and_result50[33]^and_result50[34]^and_result50[35]^and_result50[36]^and_result50[37]^and_result50[38]^and_result50[39]^and_result50[40]^and_result50[41]^and_result50[42]^and_result50[43]^and_result50[44]^and_result50[45]^and_result50[46]^and_result50[47]^and_result50[48]^and_result50[49]^and_result50[50]^and_result50[51]^and_result50[52]^and_result50[53]^and_result50[54]^and_result50[55]^and_result50[56]^and_result50[57]^and_result50[58]^and_result50[59]^and_result50[60]^and_result50[61]^and_result50[62]^and_result50[63]^and_result50[64]^and_result50[65]^and_result50[66]^and_result50[67]^and_result50[68]^and_result50[69]^and_result50[70]^and_result50[71]^and_result50[72]^and_result50[73]^and_result50[74]^and_result50[75]^and_result50[76]^and_result50[77]^and_result50[78]^and_result50[79]^and_result50[80]^and_result50[81]^and_result50[82]^and_result50[83]^and_result50[84]^and_result50[85]^and_result50[86]^and_result50[87]^and_result50[88]^and_result50[89]^and_result50[90]^and_result50[91]^and_result50[92]^and_result50[93]^and_result50[94]^and_result50[95]^and_result50[96]^and_result50[97]^and_result50[98]^and_result50[99]^and_result50[100]^and_result50[101]^and_result50[102]^and_result50[103]^and_result50[104]^and_result50[105]^and_result50[106]^and_result50[107]^and_result50[108]^and_result50[109]^and_result50[110]^and_result50[111]^and_result50[112]^and_result50[113]^and_result50[114]^and_result50[115]^and_result50[116]^and_result50[117]^and_result50[118]^and_result50[119]^and_result50[120]^and_result50[121]^and_result50[122]^and_result50[123]^and_result50[124]^and_result50[125]^and_result50[126]^and_result50[127]^and_result50[128]^and_result50[129]^and_result50[130]^and_result50[131]^and_result50[132]^and_result50[133]^and_result50[134]^and_result50[135]^and_result50[136]^and_result50[137]^and_result50[138]^and_result50[139]^and_result50[140]^and_result50[141]^and_result50[142]^and_result50[143]^and_result50[144]^and_result50[145]^and_result50[146]^and_result50[147]^and_result50[148]^and_result50[149]^and_result50[150]^and_result50[151]^and_result50[152]^and_result50[153]^and_result50[154]^and_result50[155]^and_result50[156]^and_result50[157]^and_result50[158]^and_result50[159]^and_result50[160]^and_result50[161]^and_result50[162]^and_result50[163]^and_result50[164]^and_result50[165]^and_result50[166]^and_result50[167]^and_result50[168]^and_result50[169]^and_result50[170]^and_result50[171]^and_result50[172]^and_result50[173]^and_result50[174]^and_result50[175]^and_result50[176]^and_result50[177]^and_result50[178]^and_result50[179]^and_result50[180]^and_result50[181]^and_result50[182]^and_result50[183]^and_result50[184]^and_result50[185]^and_result50[186]^and_result50[187]^and_result50[188]^and_result50[189]^and_result50[190]^and_result50[191]^and_result50[192]^and_result50[193]^and_result50[194]^and_result50[195]^and_result50[196]^and_result50[197]^and_result50[198]^and_result50[199]^and_result50[200]^and_result50[201]^and_result50[202]^and_result50[203]^and_result50[204]^and_result50[205]^and_result50[206]^and_result50[207]^and_result50[208]^and_result50[209]^and_result50[210]^and_result50[211]^and_result50[212]^and_result50[213]^and_result50[214]^and_result50[215]^and_result50[216]^and_result50[217]^and_result50[218]^and_result50[219]^and_result50[220]^and_result50[221]^and_result50[222]^and_result50[223]^and_result50[224]^and_result50[225]^and_result50[226]^and_result50[227]^and_result50[228]^and_result50[229]^and_result50[230]^and_result50[231]^and_result50[232]^and_result50[233]^and_result50[234]^and_result50[235]^and_result50[236]^and_result50[237]^and_result50[238]^and_result50[239]^and_result50[240]^and_result50[241]^and_result50[242]^and_result50[243]^and_result50[244]^and_result50[245]^and_result50[246]^and_result50[247]^and_result50[248]^and_result50[249]^and_result50[250]^and_result50[251]^and_result50[252]^and_result50[253]^and_result50[254];
assign key[51]=and_result51[0]^and_result51[1]^and_result51[2]^and_result51[3]^and_result51[4]^and_result51[5]^and_result51[6]^and_result51[7]^and_result51[8]^and_result51[9]^and_result51[10]^and_result51[11]^and_result51[12]^and_result51[13]^and_result51[14]^and_result51[15]^and_result51[16]^and_result51[17]^and_result51[18]^and_result51[19]^and_result51[20]^and_result51[21]^and_result51[22]^and_result51[23]^and_result51[24]^and_result51[25]^and_result51[26]^and_result51[27]^and_result51[28]^and_result51[29]^and_result51[30]^and_result51[31]^and_result51[32]^and_result51[33]^and_result51[34]^and_result51[35]^and_result51[36]^and_result51[37]^and_result51[38]^and_result51[39]^and_result51[40]^and_result51[41]^and_result51[42]^and_result51[43]^and_result51[44]^and_result51[45]^and_result51[46]^and_result51[47]^and_result51[48]^and_result51[49]^and_result51[50]^and_result51[51]^and_result51[52]^and_result51[53]^and_result51[54]^and_result51[55]^and_result51[56]^and_result51[57]^and_result51[58]^and_result51[59]^and_result51[60]^and_result51[61]^and_result51[62]^and_result51[63]^and_result51[64]^and_result51[65]^and_result51[66]^and_result51[67]^and_result51[68]^and_result51[69]^and_result51[70]^and_result51[71]^and_result51[72]^and_result51[73]^and_result51[74]^and_result51[75]^and_result51[76]^and_result51[77]^and_result51[78]^and_result51[79]^and_result51[80]^and_result51[81]^and_result51[82]^and_result51[83]^and_result51[84]^and_result51[85]^and_result51[86]^and_result51[87]^and_result51[88]^and_result51[89]^and_result51[90]^and_result51[91]^and_result51[92]^and_result51[93]^and_result51[94]^and_result51[95]^and_result51[96]^and_result51[97]^and_result51[98]^and_result51[99]^and_result51[100]^and_result51[101]^and_result51[102]^and_result51[103]^and_result51[104]^and_result51[105]^and_result51[106]^and_result51[107]^and_result51[108]^and_result51[109]^and_result51[110]^and_result51[111]^and_result51[112]^and_result51[113]^and_result51[114]^and_result51[115]^and_result51[116]^and_result51[117]^and_result51[118]^and_result51[119]^and_result51[120]^and_result51[121]^and_result51[122]^and_result51[123]^and_result51[124]^and_result51[125]^and_result51[126]^and_result51[127]^and_result51[128]^and_result51[129]^and_result51[130]^and_result51[131]^and_result51[132]^and_result51[133]^and_result51[134]^and_result51[135]^and_result51[136]^and_result51[137]^and_result51[138]^and_result51[139]^and_result51[140]^and_result51[141]^and_result51[142]^and_result51[143]^and_result51[144]^and_result51[145]^and_result51[146]^and_result51[147]^and_result51[148]^and_result51[149]^and_result51[150]^and_result51[151]^and_result51[152]^and_result51[153]^and_result51[154]^and_result51[155]^and_result51[156]^and_result51[157]^and_result51[158]^and_result51[159]^and_result51[160]^and_result51[161]^and_result51[162]^and_result51[163]^and_result51[164]^and_result51[165]^and_result51[166]^and_result51[167]^and_result51[168]^and_result51[169]^and_result51[170]^and_result51[171]^and_result51[172]^and_result51[173]^and_result51[174]^and_result51[175]^and_result51[176]^and_result51[177]^and_result51[178]^and_result51[179]^and_result51[180]^and_result51[181]^and_result51[182]^and_result51[183]^and_result51[184]^and_result51[185]^and_result51[186]^and_result51[187]^and_result51[188]^and_result51[189]^and_result51[190]^and_result51[191]^and_result51[192]^and_result51[193]^and_result51[194]^and_result51[195]^and_result51[196]^and_result51[197]^and_result51[198]^and_result51[199]^and_result51[200]^and_result51[201]^and_result51[202]^and_result51[203]^and_result51[204]^and_result51[205]^and_result51[206]^and_result51[207]^and_result51[208]^and_result51[209]^and_result51[210]^and_result51[211]^and_result51[212]^and_result51[213]^and_result51[214]^and_result51[215]^and_result51[216]^and_result51[217]^and_result51[218]^and_result51[219]^and_result51[220]^and_result51[221]^and_result51[222]^and_result51[223]^and_result51[224]^and_result51[225]^and_result51[226]^and_result51[227]^and_result51[228]^and_result51[229]^and_result51[230]^and_result51[231]^and_result51[232]^and_result51[233]^and_result51[234]^and_result51[235]^and_result51[236]^and_result51[237]^and_result51[238]^and_result51[239]^and_result51[240]^and_result51[241]^and_result51[242]^and_result51[243]^and_result51[244]^and_result51[245]^and_result51[246]^and_result51[247]^and_result51[248]^and_result51[249]^and_result51[250]^and_result51[251]^and_result51[252]^and_result51[253]^and_result51[254];
assign key[52]=and_result52[0]^and_result52[1]^and_result52[2]^and_result52[3]^and_result52[4]^and_result52[5]^and_result52[6]^and_result52[7]^and_result52[8]^and_result52[9]^and_result52[10]^and_result52[11]^and_result52[12]^and_result52[13]^and_result52[14]^and_result52[15]^and_result52[16]^and_result52[17]^and_result52[18]^and_result52[19]^and_result52[20]^and_result52[21]^and_result52[22]^and_result52[23]^and_result52[24]^and_result52[25]^and_result52[26]^and_result52[27]^and_result52[28]^and_result52[29]^and_result52[30]^and_result52[31]^and_result52[32]^and_result52[33]^and_result52[34]^and_result52[35]^and_result52[36]^and_result52[37]^and_result52[38]^and_result52[39]^and_result52[40]^and_result52[41]^and_result52[42]^and_result52[43]^and_result52[44]^and_result52[45]^and_result52[46]^and_result52[47]^and_result52[48]^and_result52[49]^and_result52[50]^and_result52[51]^and_result52[52]^and_result52[53]^and_result52[54]^and_result52[55]^and_result52[56]^and_result52[57]^and_result52[58]^and_result52[59]^and_result52[60]^and_result52[61]^and_result52[62]^and_result52[63]^and_result52[64]^and_result52[65]^and_result52[66]^and_result52[67]^and_result52[68]^and_result52[69]^and_result52[70]^and_result52[71]^and_result52[72]^and_result52[73]^and_result52[74]^and_result52[75]^and_result52[76]^and_result52[77]^and_result52[78]^and_result52[79]^and_result52[80]^and_result52[81]^and_result52[82]^and_result52[83]^and_result52[84]^and_result52[85]^and_result52[86]^and_result52[87]^and_result52[88]^and_result52[89]^and_result52[90]^and_result52[91]^and_result52[92]^and_result52[93]^and_result52[94]^and_result52[95]^and_result52[96]^and_result52[97]^and_result52[98]^and_result52[99]^and_result52[100]^and_result52[101]^and_result52[102]^and_result52[103]^and_result52[104]^and_result52[105]^and_result52[106]^and_result52[107]^and_result52[108]^and_result52[109]^and_result52[110]^and_result52[111]^and_result52[112]^and_result52[113]^and_result52[114]^and_result52[115]^and_result52[116]^and_result52[117]^and_result52[118]^and_result52[119]^and_result52[120]^and_result52[121]^and_result52[122]^and_result52[123]^and_result52[124]^and_result52[125]^and_result52[126]^and_result52[127]^and_result52[128]^and_result52[129]^and_result52[130]^and_result52[131]^and_result52[132]^and_result52[133]^and_result52[134]^and_result52[135]^and_result52[136]^and_result52[137]^and_result52[138]^and_result52[139]^and_result52[140]^and_result52[141]^and_result52[142]^and_result52[143]^and_result52[144]^and_result52[145]^and_result52[146]^and_result52[147]^and_result52[148]^and_result52[149]^and_result52[150]^and_result52[151]^and_result52[152]^and_result52[153]^and_result52[154]^and_result52[155]^and_result52[156]^and_result52[157]^and_result52[158]^and_result52[159]^and_result52[160]^and_result52[161]^and_result52[162]^and_result52[163]^and_result52[164]^and_result52[165]^and_result52[166]^and_result52[167]^and_result52[168]^and_result52[169]^and_result52[170]^and_result52[171]^and_result52[172]^and_result52[173]^and_result52[174]^and_result52[175]^and_result52[176]^and_result52[177]^and_result52[178]^and_result52[179]^and_result52[180]^and_result52[181]^and_result52[182]^and_result52[183]^and_result52[184]^and_result52[185]^and_result52[186]^and_result52[187]^and_result52[188]^and_result52[189]^and_result52[190]^and_result52[191]^and_result52[192]^and_result52[193]^and_result52[194]^and_result52[195]^and_result52[196]^and_result52[197]^and_result52[198]^and_result52[199]^and_result52[200]^and_result52[201]^and_result52[202]^and_result52[203]^and_result52[204]^and_result52[205]^and_result52[206]^and_result52[207]^and_result52[208]^and_result52[209]^and_result52[210]^and_result52[211]^and_result52[212]^and_result52[213]^and_result52[214]^and_result52[215]^and_result52[216]^and_result52[217]^and_result52[218]^and_result52[219]^and_result52[220]^and_result52[221]^and_result52[222]^and_result52[223]^and_result52[224]^and_result52[225]^and_result52[226]^and_result52[227]^and_result52[228]^and_result52[229]^and_result52[230]^and_result52[231]^and_result52[232]^and_result52[233]^and_result52[234]^and_result52[235]^and_result52[236]^and_result52[237]^and_result52[238]^and_result52[239]^and_result52[240]^and_result52[241]^and_result52[242]^and_result52[243]^and_result52[244]^and_result52[245]^and_result52[246]^and_result52[247]^and_result52[248]^and_result52[249]^and_result52[250]^and_result52[251]^and_result52[252]^and_result52[253]^and_result52[254];
assign key[53]=and_result53[0]^and_result53[1]^and_result53[2]^and_result53[3]^and_result53[4]^and_result53[5]^and_result53[6]^and_result53[7]^and_result53[8]^and_result53[9]^and_result53[10]^and_result53[11]^and_result53[12]^and_result53[13]^and_result53[14]^and_result53[15]^and_result53[16]^and_result53[17]^and_result53[18]^and_result53[19]^and_result53[20]^and_result53[21]^and_result53[22]^and_result53[23]^and_result53[24]^and_result53[25]^and_result53[26]^and_result53[27]^and_result53[28]^and_result53[29]^and_result53[30]^and_result53[31]^and_result53[32]^and_result53[33]^and_result53[34]^and_result53[35]^and_result53[36]^and_result53[37]^and_result53[38]^and_result53[39]^and_result53[40]^and_result53[41]^and_result53[42]^and_result53[43]^and_result53[44]^and_result53[45]^and_result53[46]^and_result53[47]^and_result53[48]^and_result53[49]^and_result53[50]^and_result53[51]^and_result53[52]^and_result53[53]^and_result53[54]^and_result53[55]^and_result53[56]^and_result53[57]^and_result53[58]^and_result53[59]^and_result53[60]^and_result53[61]^and_result53[62]^and_result53[63]^and_result53[64]^and_result53[65]^and_result53[66]^and_result53[67]^and_result53[68]^and_result53[69]^and_result53[70]^and_result53[71]^and_result53[72]^and_result53[73]^and_result53[74]^and_result53[75]^and_result53[76]^and_result53[77]^and_result53[78]^and_result53[79]^and_result53[80]^and_result53[81]^and_result53[82]^and_result53[83]^and_result53[84]^and_result53[85]^and_result53[86]^and_result53[87]^and_result53[88]^and_result53[89]^and_result53[90]^and_result53[91]^and_result53[92]^and_result53[93]^and_result53[94]^and_result53[95]^and_result53[96]^and_result53[97]^and_result53[98]^and_result53[99]^and_result53[100]^and_result53[101]^and_result53[102]^and_result53[103]^and_result53[104]^and_result53[105]^and_result53[106]^and_result53[107]^and_result53[108]^and_result53[109]^and_result53[110]^and_result53[111]^and_result53[112]^and_result53[113]^and_result53[114]^and_result53[115]^and_result53[116]^and_result53[117]^and_result53[118]^and_result53[119]^and_result53[120]^and_result53[121]^and_result53[122]^and_result53[123]^and_result53[124]^and_result53[125]^and_result53[126]^and_result53[127]^and_result53[128]^and_result53[129]^and_result53[130]^and_result53[131]^and_result53[132]^and_result53[133]^and_result53[134]^and_result53[135]^and_result53[136]^and_result53[137]^and_result53[138]^and_result53[139]^and_result53[140]^and_result53[141]^and_result53[142]^and_result53[143]^and_result53[144]^and_result53[145]^and_result53[146]^and_result53[147]^and_result53[148]^and_result53[149]^and_result53[150]^and_result53[151]^and_result53[152]^and_result53[153]^and_result53[154]^and_result53[155]^and_result53[156]^and_result53[157]^and_result53[158]^and_result53[159]^and_result53[160]^and_result53[161]^and_result53[162]^and_result53[163]^and_result53[164]^and_result53[165]^and_result53[166]^and_result53[167]^and_result53[168]^and_result53[169]^and_result53[170]^and_result53[171]^and_result53[172]^and_result53[173]^and_result53[174]^and_result53[175]^and_result53[176]^and_result53[177]^and_result53[178]^and_result53[179]^and_result53[180]^and_result53[181]^and_result53[182]^and_result53[183]^and_result53[184]^and_result53[185]^and_result53[186]^and_result53[187]^and_result53[188]^and_result53[189]^and_result53[190]^and_result53[191]^and_result53[192]^and_result53[193]^and_result53[194]^and_result53[195]^and_result53[196]^and_result53[197]^and_result53[198]^and_result53[199]^and_result53[200]^and_result53[201]^and_result53[202]^and_result53[203]^and_result53[204]^and_result53[205]^and_result53[206]^and_result53[207]^and_result53[208]^and_result53[209]^and_result53[210]^and_result53[211]^and_result53[212]^and_result53[213]^and_result53[214]^and_result53[215]^and_result53[216]^and_result53[217]^and_result53[218]^and_result53[219]^and_result53[220]^and_result53[221]^and_result53[222]^and_result53[223]^and_result53[224]^and_result53[225]^and_result53[226]^and_result53[227]^and_result53[228]^and_result53[229]^and_result53[230]^and_result53[231]^and_result53[232]^and_result53[233]^and_result53[234]^and_result53[235]^and_result53[236]^and_result53[237]^and_result53[238]^and_result53[239]^and_result53[240]^and_result53[241]^and_result53[242]^and_result53[243]^and_result53[244]^and_result53[245]^and_result53[246]^and_result53[247]^and_result53[248]^and_result53[249]^and_result53[250]^and_result53[251]^and_result53[252]^and_result53[253]^and_result53[254];
assign key[54]=and_result54[0]^and_result54[1]^and_result54[2]^and_result54[3]^and_result54[4]^and_result54[5]^and_result54[6]^and_result54[7]^and_result54[8]^and_result54[9]^and_result54[10]^and_result54[11]^and_result54[12]^and_result54[13]^and_result54[14]^and_result54[15]^and_result54[16]^and_result54[17]^and_result54[18]^and_result54[19]^and_result54[20]^and_result54[21]^and_result54[22]^and_result54[23]^and_result54[24]^and_result54[25]^and_result54[26]^and_result54[27]^and_result54[28]^and_result54[29]^and_result54[30]^and_result54[31]^and_result54[32]^and_result54[33]^and_result54[34]^and_result54[35]^and_result54[36]^and_result54[37]^and_result54[38]^and_result54[39]^and_result54[40]^and_result54[41]^and_result54[42]^and_result54[43]^and_result54[44]^and_result54[45]^and_result54[46]^and_result54[47]^and_result54[48]^and_result54[49]^and_result54[50]^and_result54[51]^and_result54[52]^and_result54[53]^and_result54[54]^and_result54[55]^and_result54[56]^and_result54[57]^and_result54[58]^and_result54[59]^and_result54[60]^and_result54[61]^and_result54[62]^and_result54[63]^and_result54[64]^and_result54[65]^and_result54[66]^and_result54[67]^and_result54[68]^and_result54[69]^and_result54[70]^and_result54[71]^and_result54[72]^and_result54[73]^and_result54[74]^and_result54[75]^and_result54[76]^and_result54[77]^and_result54[78]^and_result54[79]^and_result54[80]^and_result54[81]^and_result54[82]^and_result54[83]^and_result54[84]^and_result54[85]^and_result54[86]^and_result54[87]^and_result54[88]^and_result54[89]^and_result54[90]^and_result54[91]^and_result54[92]^and_result54[93]^and_result54[94]^and_result54[95]^and_result54[96]^and_result54[97]^and_result54[98]^and_result54[99]^and_result54[100]^and_result54[101]^and_result54[102]^and_result54[103]^and_result54[104]^and_result54[105]^and_result54[106]^and_result54[107]^and_result54[108]^and_result54[109]^and_result54[110]^and_result54[111]^and_result54[112]^and_result54[113]^and_result54[114]^and_result54[115]^and_result54[116]^and_result54[117]^and_result54[118]^and_result54[119]^and_result54[120]^and_result54[121]^and_result54[122]^and_result54[123]^and_result54[124]^and_result54[125]^and_result54[126]^and_result54[127]^and_result54[128]^and_result54[129]^and_result54[130]^and_result54[131]^and_result54[132]^and_result54[133]^and_result54[134]^and_result54[135]^and_result54[136]^and_result54[137]^and_result54[138]^and_result54[139]^and_result54[140]^and_result54[141]^and_result54[142]^and_result54[143]^and_result54[144]^and_result54[145]^and_result54[146]^and_result54[147]^and_result54[148]^and_result54[149]^and_result54[150]^and_result54[151]^and_result54[152]^and_result54[153]^and_result54[154]^and_result54[155]^and_result54[156]^and_result54[157]^and_result54[158]^and_result54[159]^and_result54[160]^and_result54[161]^and_result54[162]^and_result54[163]^and_result54[164]^and_result54[165]^and_result54[166]^and_result54[167]^and_result54[168]^and_result54[169]^and_result54[170]^and_result54[171]^and_result54[172]^and_result54[173]^and_result54[174]^and_result54[175]^and_result54[176]^and_result54[177]^and_result54[178]^and_result54[179]^and_result54[180]^and_result54[181]^and_result54[182]^and_result54[183]^and_result54[184]^and_result54[185]^and_result54[186]^and_result54[187]^and_result54[188]^and_result54[189]^and_result54[190]^and_result54[191]^and_result54[192]^and_result54[193]^and_result54[194]^and_result54[195]^and_result54[196]^and_result54[197]^and_result54[198]^and_result54[199]^and_result54[200]^and_result54[201]^and_result54[202]^and_result54[203]^and_result54[204]^and_result54[205]^and_result54[206]^and_result54[207]^and_result54[208]^and_result54[209]^and_result54[210]^and_result54[211]^and_result54[212]^and_result54[213]^and_result54[214]^and_result54[215]^and_result54[216]^and_result54[217]^and_result54[218]^and_result54[219]^and_result54[220]^and_result54[221]^and_result54[222]^and_result54[223]^and_result54[224]^and_result54[225]^and_result54[226]^and_result54[227]^and_result54[228]^and_result54[229]^and_result54[230]^and_result54[231]^and_result54[232]^and_result54[233]^and_result54[234]^and_result54[235]^and_result54[236]^and_result54[237]^and_result54[238]^and_result54[239]^and_result54[240]^and_result54[241]^and_result54[242]^and_result54[243]^and_result54[244]^and_result54[245]^and_result54[246]^and_result54[247]^and_result54[248]^and_result54[249]^and_result54[250]^and_result54[251]^and_result54[252]^and_result54[253]^and_result54[254];
assign key[55]=and_result55[0]^and_result55[1]^and_result55[2]^and_result55[3]^and_result55[4]^and_result55[5]^and_result55[6]^and_result55[7]^and_result55[8]^and_result55[9]^and_result55[10]^and_result55[11]^and_result55[12]^and_result55[13]^and_result55[14]^and_result55[15]^and_result55[16]^and_result55[17]^and_result55[18]^and_result55[19]^and_result55[20]^and_result55[21]^and_result55[22]^and_result55[23]^and_result55[24]^and_result55[25]^and_result55[26]^and_result55[27]^and_result55[28]^and_result55[29]^and_result55[30]^and_result55[31]^and_result55[32]^and_result55[33]^and_result55[34]^and_result55[35]^and_result55[36]^and_result55[37]^and_result55[38]^and_result55[39]^and_result55[40]^and_result55[41]^and_result55[42]^and_result55[43]^and_result55[44]^and_result55[45]^and_result55[46]^and_result55[47]^and_result55[48]^and_result55[49]^and_result55[50]^and_result55[51]^and_result55[52]^and_result55[53]^and_result55[54]^and_result55[55]^and_result55[56]^and_result55[57]^and_result55[58]^and_result55[59]^and_result55[60]^and_result55[61]^and_result55[62]^and_result55[63]^and_result55[64]^and_result55[65]^and_result55[66]^and_result55[67]^and_result55[68]^and_result55[69]^and_result55[70]^and_result55[71]^and_result55[72]^and_result55[73]^and_result55[74]^and_result55[75]^and_result55[76]^and_result55[77]^and_result55[78]^and_result55[79]^and_result55[80]^and_result55[81]^and_result55[82]^and_result55[83]^and_result55[84]^and_result55[85]^and_result55[86]^and_result55[87]^and_result55[88]^and_result55[89]^and_result55[90]^and_result55[91]^and_result55[92]^and_result55[93]^and_result55[94]^and_result55[95]^and_result55[96]^and_result55[97]^and_result55[98]^and_result55[99]^and_result55[100]^and_result55[101]^and_result55[102]^and_result55[103]^and_result55[104]^and_result55[105]^and_result55[106]^and_result55[107]^and_result55[108]^and_result55[109]^and_result55[110]^and_result55[111]^and_result55[112]^and_result55[113]^and_result55[114]^and_result55[115]^and_result55[116]^and_result55[117]^and_result55[118]^and_result55[119]^and_result55[120]^and_result55[121]^and_result55[122]^and_result55[123]^and_result55[124]^and_result55[125]^and_result55[126]^and_result55[127]^and_result55[128]^and_result55[129]^and_result55[130]^and_result55[131]^and_result55[132]^and_result55[133]^and_result55[134]^and_result55[135]^and_result55[136]^and_result55[137]^and_result55[138]^and_result55[139]^and_result55[140]^and_result55[141]^and_result55[142]^and_result55[143]^and_result55[144]^and_result55[145]^and_result55[146]^and_result55[147]^and_result55[148]^and_result55[149]^and_result55[150]^and_result55[151]^and_result55[152]^and_result55[153]^and_result55[154]^and_result55[155]^and_result55[156]^and_result55[157]^and_result55[158]^and_result55[159]^and_result55[160]^and_result55[161]^and_result55[162]^and_result55[163]^and_result55[164]^and_result55[165]^and_result55[166]^and_result55[167]^and_result55[168]^and_result55[169]^and_result55[170]^and_result55[171]^and_result55[172]^and_result55[173]^and_result55[174]^and_result55[175]^and_result55[176]^and_result55[177]^and_result55[178]^and_result55[179]^and_result55[180]^and_result55[181]^and_result55[182]^and_result55[183]^and_result55[184]^and_result55[185]^and_result55[186]^and_result55[187]^and_result55[188]^and_result55[189]^and_result55[190]^and_result55[191]^and_result55[192]^and_result55[193]^and_result55[194]^and_result55[195]^and_result55[196]^and_result55[197]^and_result55[198]^and_result55[199]^and_result55[200]^and_result55[201]^and_result55[202]^and_result55[203]^and_result55[204]^and_result55[205]^and_result55[206]^and_result55[207]^and_result55[208]^and_result55[209]^and_result55[210]^and_result55[211]^and_result55[212]^and_result55[213]^and_result55[214]^and_result55[215]^and_result55[216]^and_result55[217]^and_result55[218]^and_result55[219]^and_result55[220]^and_result55[221]^and_result55[222]^and_result55[223]^and_result55[224]^and_result55[225]^and_result55[226]^and_result55[227]^and_result55[228]^and_result55[229]^and_result55[230]^and_result55[231]^and_result55[232]^and_result55[233]^and_result55[234]^and_result55[235]^and_result55[236]^and_result55[237]^and_result55[238]^and_result55[239]^and_result55[240]^and_result55[241]^and_result55[242]^and_result55[243]^and_result55[244]^and_result55[245]^and_result55[246]^and_result55[247]^and_result55[248]^and_result55[249]^and_result55[250]^and_result55[251]^and_result55[252]^and_result55[253]^and_result55[254];
assign key[56]=and_result56[0]^and_result56[1]^and_result56[2]^and_result56[3]^and_result56[4]^and_result56[5]^and_result56[6]^and_result56[7]^and_result56[8]^and_result56[9]^and_result56[10]^and_result56[11]^and_result56[12]^and_result56[13]^and_result56[14]^and_result56[15]^and_result56[16]^and_result56[17]^and_result56[18]^and_result56[19]^and_result56[20]^and_result56[21]^and_result56[22]^and_result56[23]^and_result56[24]^and_result56[25]^and_result56[26]^and_result56[27]^and_result56[28]^and_result56[29]^and_result56[30]^and_result56[31]^and_result56[32]^and_result56[33]^and_result56[34]^and_result56[35]^and_result56[36]^and_result56[37]^and_result56[38]^and_result56[39]^and_result56[40]^and_result56[41]^and_result56[42]^and_result56[43]^and_result56[44]^and_result56[45]^and_result56[46]^and_result56[47]^and_result56[48]^and_result56[49]^and_result56[50]^and_result56[51]^and_result56[52]^and_result56[53]^and_result56[54]^and_result56[55]^and_result56[56]^and_result56[57]^and_result56[58]^and_result56[59]^and_result56[60]^and_result56[61]^and_result56[62]^and_result56[63]^and_result56[64]^and_result56[65]^and_result56[66]^and_result56[67]^and_result56[68]^and_result56[69]^and_result56[70]^and_result56[71]^and_result56[72]^and_result56[73]^and_result56[74]^and_result56[75]^and_result56[76]^and_result56[77]^and_result56[78]^and_result56[79]^and_result56[80]^and_result56[81]^and_result56[82]^and_result56[83]^and_result56[84]^and_result56[85]^and_result56[86]^and_result56[87]^and_result56[88]^and_result56[89]^and_result56[90]^and_result56[91]^and_result56[92]^and_result56[93]^and_result56[94]^and_result56[95]^and_result56[96]^and_result56[97]^and_result56[98]^and_result56[99]^and_result56[100]^and_result56[101]^and_result56[102]^and_result56[103]^and_result56[104]^and_result56[105]^and_result56[106]^and_result56[107]^and_result56[108]^and_result56[109]^and_result56[110]^and_result56[111]^and_result56[112]^and_result56[113]^and_result56[114]^and_result56[115]^and_result56[116]^and_result56[117]^and_result56[118]^and_result56[119]^and_result56[120]^and_result56[121]^and_result56[122]^and_result56[123]^and_result56[124]^and_result56[125]^and_result56[126]^and_result56[127]^and_result56[128]^and_result56[129]^and_result56[130]^and_result56[131]^and_result56[132]^and_result56[133]^and_result56[134]^and_result56[135]^and_result56[136]^and_result56[137]^and_result56[138]^and_result56[139]^and_result56[140]^and_result56[141]^and_result56[142]^and_result56[143]^and_result56[144]^and_result56[145]^and_result56[146]^and_result56[147]^and_result56[148]^and_result56[149]^and_result56[150]^and_result56[151]^and_result56[152]^and_result56[153]^and_result56[154]^and_result56[155]^and_result56[156]^and_result56[157]^and_result56[158]^and_result56[159]^and_result56[160]^and_result56[161]^and_result56[162]^and_result56[163]^and_result56[164]^and_result56[165]^and_result56[166]^and_result56[167]^and_result56[168]^and_result56[169]^and_result56[170]^and_result56[171]^and_result56[172]^and_result56[173]^and_result56[174]^and_result56[175]^and_result56[176]^and_result56[177]^and_result56[178]^and_result56[179]^and_result56[180]^and_result56[181]^and_result56[182]^and_result56[183]^and_result56[184]^and_result56[185]^and_result56[186]^and_result56[187]^and_result56[188]^and_result56[189]^and_result56[190]^and_result56[191]^and_result56[192]^and_result56[193]^and_result56[194]^and_result56[195]^and_result56[196]^and_result56[197]^and_result56[198]^and_result56[199]^and_result56[200]^and_result56[201]^and_result56[202]^and_result56[203]^and_result56[204]^and_result56[205]^and_result56[206]^and_result56[207]^and_result56[208]^and_result56[209]^and_result56[210]^and_result56[211]^and_result56[212]^and_result56[213]^and_result56[214]^and_result56[215]^and_result56[216]^and_result56[217]^and_result56[218]^and_result56[219]^and_result56[220]^and_result56[221]^and_result56[222]^and_result56[223]^and_result56[224]^and_result56[225]^and_result56[226]^and_result56[227]^and_result56[228]^and_result56[229]^and_result56[230]^and_result56[231]^and_result56[232]^and_result56[233]^and_result56[234]^and_result56[235]^and_result56[236]^and_result56[237]^and_result56[238]^and_result56[239]^and_result56[240]^and_result56[241]^and_result56[242]^and_result56[243]^and_result56[244]^and_result56[245]^and_result56[246]^and_result56[247]^and_result56[248]^and_result56[249]^and_result56[250]^and_result56[251]^and_result56[252]^and_result56[253]^and_result56[254];
assign key[57]=and_result57[0]^and_result57[1]^and_result57[2]^and_result57[3]^and_result57[4]^and_result57[5]^and_result57[6]^and_result57[7]^and_result57[8]^and_result57[9]^and_result57[10]^and_result57[11]^and_result57[12]^and_result57[13]^and_result57[14]^and_result57[15]^and_result57[16]^and_result57[17]^and_result57[18]^and_result57[19]^and_result57[20]^and_result57[21]^and_result57[22]^and_result57[23]^and_result57[24]^and_result57[25]^and_result57[26]^and_result57[27]^and_result57[28]^and_result57[29]^and_result57[30]^and_result57[31]^and_result57[32]^and_result57[33]^and_result57[34]^and_result57[35]^and_result57[36]^and_result57[37]^and_result57[38]^and_result57[39]^and_result57[40]^and_result57[41]^and_result57[42]^and_result57[43]^and_result57[44]^and_result57[45]^and_result57[46]^and_result57[47]^and_result57[48]^and_result57[49]^and_result57[50]^and_result57[51]^and_result57[52]^and_result57[53]^and_result57[54]^and_result57[55]^and_result57[56]^and_result57[57]^and_result57[58]^and_result57[59]^and_result57[60]^and_result57[61]^and_result57[62]^and_result57[63]^and_result57[64]^and_result57[65]^and_result57[66]^and_result57[67]^and_result57[68]^and_result57[69]^and_result57[70]^and_result57[71]^and_result57[72]^and_result57[73]^and_result57[74]^and_result57[75]^and_result57[76]^and_result57[77]^and_result57[78]^and_result57[79]^and_result57[80]^and_result57[81]^and_result57[82]^and_result57[83]^and_result57[84]^and_result57[85]^and_result57[86]^and_result57[87]^and_result57[88]^and_result57[89]^and_result57[90]^and_result57[91]^and_result57[92]^and_result57[93]^and_result57[94]^and_result57[95]^and_result57[96]^and_result57[97]^and_result57[98]^and_result57[99]^and_result57[100]^and_result57[101]^and_result57[102]^and_result57[103]^and_result57[104]^and_result57[105]^and_result57[106]^and_result57[107]^and_result57[108]^and_result57[109]^and_result57[110]^and_result57[111]^and_result57[112]^and_result57[113]^and_result57[114]^and_result57[115]^and_result57[116]^and_result57[117]^and_result57[118]^and_result57[119]^and_result57[120]^and_result57[121]^and_result57[122]^and_result57[123]^and_result57[124]^and_result57[125]^and_result57[126]^and_result57[127]^and_result57[128]^and_result57[129]^and_result57[130]^and_result57[131]^and_result57[132]^and_result57[133]^and_result57[134]^and_result57[135]^and_result57[136]^and_result57[137]^and_result57[138]^and_result57[139]^and_result57[140]^and_result57[141]^and_result57[142]^and_result57[143]^and_result57[144]^and_result57[145]^and_result57[146]^and_result57[147]^and_result57[148]^and_result57[149]^and_result57[150]^and_result57[151]^and_result57[152]^and_result57[153]^and_result57[154]^and_result57[155]^and_result57[156]^and_result57[157]^and_result57[158]^and_result57[159]^and_result57[160]^and_result57[161]^and_result57[162]^and_result57[163]^and_result57[164]^and_result57[165]^and_result57[166]^and_result57[167]^and_result57[168]^and_result57[169]^and_result57[170]^and_result57[171]^and_result57[172]^and_result57[173]^and_result57[174]^and_result57[175]^and_result57[176]^and_result57[177]^and_result57[178]^and_result57[179]^and_result57[180]^and_result57[181]^and_result57[182]^and_result57[183]^and_result57[184]^and_result57[185]^and_result57[186]^and_result57[187]^and_result57[188]^and_result57[189]^and_result57[190]^and_result57[191]^and_result57[192]^and_result57[193]^and_result57[194]^and_result57[195]^and_result57[196]^and_result57[197]^and_result57[198]^and_result57[199]^and_result57[200]^and_result57[201]^and_result57[202]^and_result57[203]^and_result57[204]^and_result57[205]^and_result57[206]^and_result57[207]^and_result57[208]^and_result57[209]^and_result57[210]^and_result57[211]^and_result57[212]^and_result57[213]^and_result57[214]^and_result57[215]^and_result57[216]^and_result57[217]^and_result57[218]^and_result57[219]^and_result57[220]^and_result57[221]^and_result57[222]^and_result57[223]^and_result57[224]^and_result57[225]^and_result57[226]^and_result57[227]^and_result57[228]^and_result57[229]^and_result57[230]^and_result57[231]^and_result57[232]^and_result57[233]^and_result57[234]^and_result57[235]^and_result57[236]^and_result57[237]^and_result57[238]^and_result57[239]^and_result57[240]^and_result57[241]^and_result57[242]^and_result57[243]^and_result57[244]^and_result57[245]^and_result57[246]^and_result57[247]^and_result57[248]^and_result57[249]^and_result57[250]^and_result57[251]^and_result57[252]^and_result57[253]^and_result57[254];
assign key[58]=and_result58[0]^and_result58[1]^and_result58[2]^and_result58[3]^and_result58[4]^and_result58[5]^and_result58[6]^and_result58[7]^and_result58[8]^and_result58[9]^and_result58[10]^and_result58[11]^and_result58[12]^and_result58[13]^and_result58[14]^and_result58[15]^and_result58[16]^and_result58[17]^and_result58[18]^and_result58[19]^and_result58[20]^and_result58[21]^and_result58[22]^and_result58[23]^and_result58[24]^and_result58[25]^and_result58[26]^and_result58[27]^and_result58[28]^and_result58[29]^and_result58[30]^and_result58[31]^and_result58[32]^and_result58[33]^and_result58[34]^and_result58[35]^and_result58[36]^and_result58[37]^and_result58[38]^and_result58[39]^and_result58[40]^and_result58[41]^and_result58[42]^and_result58[43]^and_result58[44]^and_result58[45]^and_result58[46]^and_result58[47]^and_result58[48]^and_result58[49]^and_result58[50]^and_result58[51]^and_result58[52]^and_result58[53]^and_result58[54]^and_result58[55]^and_result58[56]^and_result58[57]^and_result58[58]^and_result58[59]^and_result58[60]^and_result58[61]^and_result58[62]^and_result58[63]^and_result58[64]^and_result58[65]^and_result58[66]^and_result58[67]^and_result58[68]^and_result58[69]^and_result58[70]^and_result58[71]^and_result58[72]^and_result58[73]^and_result58[74]^and_result58[75]^and_result58[76]^and_result58[77]^and_result58[78]^and_result58[79]^and_result58[80]^and_result58[81]^and_result58[82]^and_result58[83]^and_result58[84]^and_result58[85]^and_result58[86]^and_result58[87]^and_result58[88]^and_result58[89]^and_result58[90]^and_result58[91]^and_result58[92]^and_result58[93]^and_result58[94]^and_result58[95]^and_result58[96]^and_result58[97]^and_result58[98]^and_result58[99]^and_result58[100]^and_result58[101]^and_result58[102]^and_result58[103]^and_result58[104]^and_result58[105]^and_result58[106]^and_result58[107]^and_result58[108]^and_result58[109]^and_result58[110]^and_result58[111]^and_result58[112]^and_result58[113]^and_result58[114]^and_result58[115]^and_result58[116]^and_result58[117]^and_result58[118]^and_result58[119]^and_result58[120]^and_result58[121]^and_result58[122]^and_result58[123]^and_result58[124]^and_result58[125]^and_result58[126]^and_result58[127]^and_result58[128]^and_result58[129]^and_result58[130]^and_result58[131]^and_result58[132]^and_result58[133]^and_result58[134]^and_result58[135]^and_result58[136]^and_result58[137]^and_result58[138]^and_result58[139]^and_result58[140]^and_result58[141]^and_result58[142]^and_result58[143]^and_result58[144]^and_result58[145]^and_result58[146]^and_result58[147]^and_result58[148]^and_result58[149]^and_result58[150]^and_result58[151]^and_result58[152]^and_result58[153]^and_result58[154]^and_result58[155]^and_result58[156]^and_result58[157]^and_result58[158]^and_result58[159]^and_result58[160]^and_result58[161]^and_result58[162]^and_result58[163]^and_result58[164]^and_result58[165]^and_result58[166]^and_result58[167]^and_result58[168]^and_result58[169]^and_result58[170]^and_result58[171]^and_result58[172]^and_result58[173]^and_result58[174]^and_result58[175]^and_result58[176]^and_result58[177]^and_result58[178]^and_result58[179]^and_result58[180]^and_result58[181]^and_result58[182]^and_result58[183]^and_result58[184]^and_result58[185]^and_result58[186]^and_result58[187]^and_result58[188]^and_result58[189]^and_result58[190]^and_result58[191]^and_result58[192]^and_result58[193]^and_result58[194]^and_result58[195]^and_result58[196]^and_result58[197]^and_result58[198]^and_result58[199]^and_result58[200]^and_result58[201]^and_result58[202]^and_result58[203]^and_result58[204]^and_result58[205]^and_result58[206]^and_result58[207]^and_result58[208]^and_result58[209]^and_result58[210]^and_result58[211]^and_result58[212]^and_result58[213]^and_result58[214]^and_result58[215]^and_result58[216]^and_result58[217]^and_result58[218]^and_result58[219]^and_result58[220]^and_result58[221]^and_result58[222]^and_result58[223]^and_result58[224]^and_result58[225]^and_result58[226]^and_result58[227]^and_result58[228]^and_result58[229]^and_result58[230]^and_result58[231]^and_result58[232]^and_result58[233]^and_result58[234]^and_result58[235]^and_result58[236]^and_result58[237]^and_result58[238]^and_result58[239]^and_result58[240]^and_result58[241]^and_result58[242]^and_result58[243]^and_result58[244]^and_result58[245]^and_result58[246]^and_result58[247]^and_result58[248]^and_result58[249]^and_result58[250]^and_result58[251]^and_result58[252]^and_result58[253]^and_result58[254];
assign key[59]=and_result59[0]^and_result59[1]^and_result59[2]^and_result59[3]^and_result59[4]^and_result59[5]^and_result59[6]^and_result59[7]^and_result59[8]^and_result59[9]^and_result59[10]^and_result59[11]^and_result59[12]^and_result59[13]^and_result59[14]^and_result59[15]^and_result59[16]^and_result59[17]^and_result59[18]^and_result59[19]^and_result59[20]^and_result59[21]^and_result59[22]^and_result59[23]^and_result59[24]^and_result59[25]^and_result59[26]^and_result59[27]^and_result59[28]^and_result59[29]^and_result59[30]^and_result59[31]^and_result59[32]^and_result59[33]^and_result59[34]^and_result59[35]^and_result59[36]^and_result59[37]^and_result59[38]^and_result59[39]^and_result59[40]^and_result59[41]^and_result59[42]^and_result59[43]^and_result59[44]^and_result59[45]^and_result59[46]^and_result59[47]^and_result59[48]^and_result59[49]^and_result59[50]^and_result59[51]^and_result59[52]^and_result59[53]^and_result59[54]^and_result59[55]^and_result59[56]^and_result59[57]^and_result59[58]^and_result59[59]^and_result59[60]^and_result59[61]^and_result59[62]^and_result59[63]^and_result59[64]^and_result59[65]^and_result59[66]^and_result59[67]^and_result59[68]^and_result59[69]^and_result59[70]^and_result59[71]^and_result59[72]^and_result59[73]^and_result59[74]^and_result59[75]^and_result59[76]^and_result59[77]^and_result59[78]^and_result59[79]^and_result59[80]^and_result59[81]^and_result59[82]^and_result59[83]^and_result59[84]^and_result59[85]^and_result59[86]^and_result59[87]^and_result59[88]^and_result59[89]^and_result59[90]^and_result59[91]^and_result59[92]^and_result59[93]^and_result59[94]^and_result59[95]^and_result59[96]^and_result59[97]^and_result59[98]^and_result59[99]^and_result59[100]^and_result59[101]^and_result59[102]^and_result59[103]^and_result59[104]^and_result59[105]^and_result59[106]^and_result59[107]^and_result59[108]^and_result59[109]^and_result59[110]^and_result59[111]^and_result59[112]^and_result59[113]^and_result59[114]^and_result59[115]^and_result59[116]^and_result59[117]^and_result59[118]^and_result59[119]^and_result59[120]^and_result59[121]^and_result59[122]^and_result59[123]^and_result59[124]^and_result59[125]^and_result59[126]^and_result59[127]^and_result59[128]^and_result59[129]^and_result59[130]^and_result59[131]^and_result59[132]^and_result59[133]^and_result59[134]^and_result59[135]^and_result59[136]^and_result59[137]^and_result59[138]^and_result59[139]^and_result59[140]^and_result59[141]^and_result59[142]^and_result59[143]^and_result59[144]^and_result59[145]^and_result59[146]^and_result59[147]^and_result59[148]^and_result59[149]^and_result59[150]^and_result59[151]^and_result59[152]^and_result59[153]^and_result59[154]^and_result59[155]^and_result59[156]^and_result59[157]^and_result59[158]^and_result59[159]^and_result59[160]^and_result59[161]^and_result59[162]^and_result59[163]^and_result59[164]^and_result59[165]^and_result59[166]^and_result59[167]^and_result59[168]^and_result59[169]^and_result59[170]^and_result59[171]^and_result59[172]^and_result59[173]^and_result59[174]^and_result59[175]^and_result59[176]^and_result59[177]^and_result59[178]^and_result59[179]^and_result59[180]^and_result59[181]^and_result59[182]^and_result59[183]^and_result59[184]^and_result59[185]^and_result59[186]^and_result59[187]^and_result59[188]^and_result59[189]^and_result59[190]^and_result59[191]^and_result59[192]^and_result59[193]^and_result59[194]^and_result59[195]^and_result59[196]^and_result59[197]^and_result59[198]^and_result59[199]^and_result59[200]^and_result59[201]^and_result59[202]^and_result59[203]^and_result59[204]^and_result59[205]^and_result59[206]^and_result59[207]^and_result59[208]^and_result59[209]^and_result59[210]^and_result59[211]^and_result59[212]^and_result59[213]^and_result59[214]^and_result59[215]^and_result59[216]^and_result59[217]^and_result59[218]^and_result59[219]^and_result59[220]^and_result59[221]^and_result59[222]^and_result59[223]^and_result59[224]^and_result59[225]^and_result59[226]^and_result59[227]^and_result59[228]^and_result59[229]^and_result59[230]^and_result59[231]^and_result59[232]^and_result59[233]^and_result59[234]^and_result59[235]^and_result59[236]^and_result59[237]^and_result59[238]^and_result59[239]^and_result59[240]^and_result59[241]^and_result59[242]^and_result59[243]^and_result59[244]^and_result59[245]^and_result59[246]^and_result59[247]^and_result59[248]^and_result59[249]^and_result59[250]^and_result59[251]^and_result59[252]^and_result59[253]^and_result59[254];
assign key[60]=and_result60[0]^and_result60[1]^and_result60[2]^and_result60[3]^and_result60[4]^and_result60[5]^and_result60[6]^and_result60[7]^and_result60[8]^and_result60[9]^and_result60[10]^and_result60[11]^and_result60[12]^and_result60[13]^and_result60[14]^and_result60[15]^and_result60[16]^and_result60[17]^and_result60[18]^and_result60[19]^and_result60[20]^and_result60[21]^and_result60[22]^and_result60[23]^and_result60[24]^and_result60[25]^and_result60[26]^and_result60[27]^and_result60[28]^and_result60[29]^and_result60[30]^and_result60[31]^and_result60[32]^and_result60[33]^and_result60[34]^and_result60[35]^and_result60[36]^and_result60[37]^and_result60[38]^and_result60[39]^and_result60[40]^and_result60[41]^and_result60[42]^and_result60[43]^and_result60[44]^and_result60[45]^and_result60[46]^and_result60[47]^and_result60[48]^and_result60[49]^and_result60[50]^and_result60[51]^and_result60[52]^and_result60[53]^and_result60[54]^and_result60[55]^and_result60[56]^and_result60[57]^and_result60[58]^and_result60[59]^and_result60[60]^and_result60[61]^and_result60[62]^and_result60[63]^and_result60[64]^and_result60[65]^and_result60[66]^and_result60[67]^and_result60[68]^and_result60[69]^and_result60[70]^and_result60[71]^and_result60[72]^and_result60[73]^and_result60[74]^and_result60[75]^and_result60[76]^and_result60[77]^and_result60[78]^and_result60[79]^and_result60[80]^and_result60[81]^and_result60[82]^and_result60[83]^and_result60[84]^and_result60[85]^and_result60[86]^and_result60[87]^and_result60[88]^and_result60[89]^and_result60[90]^and_result60[91]^and_result60[92]^and_result60[93]^and_result60[94]^and_result60[95]^and_result60[96]^and_result60[97]^and_result60[98]^and_result60[99]^and_result60[100]^and_result60[101]^and_result60[102]^and_result60[103]^and_result60[104]^and_result60[105]^and_result60[106]^and_result60[107]^and_result60[108]^and_result60[109]^and_result60[110]^and_result60[111]^and_result60[112]^and_result60[113]^and_result60[114]^and_result60[115]^and_result60[116]^and_result60[117]^and_result60[118]^and_result60[119]^and_result60[120]^and_result60[121]^and_result60[122]^and_result60[123]^and_result60[124]^and_result60[125]^and_result60[126]^and_result60[127]^and_result60[128]^and_result60[129]^and_result60[130]^and_result60[131]^and_result60[132]^and_result60[133]^and_result60[134]^and_result60[135]^and_result60[136]^and_result60[137]^and_result60[138]^and_result60[139]^and_result60[140]^and_result60[141]^and_result60[142]^and_result60[143]^and_result60[144]^and_result60[145]^and_result60[146]^and_result60[147]^and_result60[148]^and_result60[149]^and_result60[150]^and_result60[151]^and_result60[152]^and_result60[153]^and_result60[154]^and_result60[155]^and_result60[156]^and_result60[157]^and_result60[158]^and_result60[159]^and_result60[160]^and_result60[161]^and_result60[162]^and_result60[163]^and_result60[164]^and_result60[165]^and_result60[166]^and_result60[167]^and_result60[168]^and_result60[169]^and_result60[170]^and_result60[171]^and_result60[172]^and_result60[173]^and_result60[174]^and_result60[175]^and_result60[176]^and_result60[177]^and_result60[178]^and_result60[179]^and_result60[180]^and_result60[181]^and_result60[182]^and_result60[183]^and_result60[184]^and_result60[185]^and_result60[186]^and_result60[187]^and_result60[188]^and_result60[189]^and_result60[190]^and_result60[191]^and_result60[192]^and_result60[193]^and_result60[194]^and_result60[195]^and_result60[196]^and_result60[197]^and_result60[198]^and_result60[199]^and_result60[200]^and_result60[201]^and_result60[202]^and_result60[203]^and_result60[204]^and_result60[205]^and_result60[206]^and_result60[207]^and_result60[208]^and_result60[209]^and_result60[210]^and_result60[211]^and_result60[212]^and_result60[213]^and_result60[214]^and_result60[215]^and_result60[216]^and_result60[217]^and_result60[218]^and_result60[219]^and_result60[220]^and_result60[221]^and_result60[222]^and_result60[223]^and_result60[224]^and_result60[225]^and_result60[226]^and_result60[227]^and_result60[228]^and_result60[229]^and_result60[230]^and_result60[231]^and_result60[232]^and_result60[233]^and_result60[234]^and_result60[235]^and_result60[236]^and_result60[237]^and_result60[238]^and_result60[239]^and_result60[240]^and_result60[241]^and_result60[242]^and_result60[243]^and_result60[244]^and_result60[245]^and_result60[246]^and_result60[247]^and_result60[248]^and_result60[249]^and_result60[250]^and_result60[251]^and_result60[252]^and_result60[253]^and_result60[254];
assign key[61]=and_result61[0]^and_result61[1]^and_result61[2]^and_result61[3]^and_result61[4]^and_result61[5]^and_result61[6]^and_result61[7]^and_result61[8]^and_result61[9]^and_result61[10]^and_result61[11]^and_result61[12]^and_result61[13]^and_result61[14]^and_result61[15]^and_result61[16]^and_result61[17]^and_result61[18]^and_result61[19]^and_result61[20]^and_result61[21]^and_result61[22]^and_result61[23]^and_result61[24]^and_result61[25]^and_result61[26]^and_result61[27]^and_result61[28]^and_result61[29]^and_result61[30]^and_result61[31]^and_result61[32]^and_result61[33]^and_result61[34]^and_result61[35]^and_result61[36]^and_result61[37]^and_result61[38]^and_result61[39]^and_result61[40]^and_result61[41]^and_result61[42]^and_result61[43]^and_result61[44]^and_result61[45]^and_result61[46]^and_result61[47]^and_result61[48]^and_result61[49]^and_result61[50]^and_result61[51]^and_result61[52]^and_result61[53]^and_result61[54]^and_result61[55]^and_result61[56]^and_result61[57]^and_result61[58]^and_result61[59]^and_result61[60]^and_result61[61]^and_result61[62]^and_result61[63]^and_result61[64]^and_result61[65]^and_result61[66]^and_result61[67]^and_result61[68]^and_result61[69]^and_result61[70]^and_result61[71]^and_result61[72]^and_result61[73]^and_result61[74]^and_result61[75]^and_result61[76]^and_result61[77]^and_result61[78]^and_result61[79]^and_result61[80]^and_result61[81]^and_result61[82]^and_result61[83]^and_result61[84]^and_result61[85]^and_result61[86]^and_result61[87]^and_result61[88]^and_result61[89]^and_result61[90]^and_result61[91]^and_result61[92]^and_result61[93]^and_result61[94]^and_result61[95]^and_result61[96]^and_result61[97]^and_result61[98]^and_result61[99]^and_result61[100]^and_result61[101]^and_result61[102]^and_result61[103]^and_result61[104]^and_result61[105]^and_result61[106]^and_result61[107]^and_result61[108]^and_result61[109]^and_result61[110]^and_result61[111]^and_result61[112]^and_result61[113]^and_result61[114]^and_result61[115]^and_result61[116]^and_result61[117]^and_result61[118]^and_result61[119]^and_result61[120]^and_result61[121]^and_result61[122]^and_result61[123]^and_result61[124]^and_result61[125]^and_result61[126]^and_result61[127]^and_result61[128]^and_result61[129]^and_result61[130]^and_result61[131]^and_result61[132]^and_result61[133]^and_result61[134]^and_result61[135]^and_result61[136]^and_result61[137]^and_result61[138]^and_result61[139]^and_result61[140]^and_result61[141]^and_result61[142]^and_result61[143]^and_result61[144]^and_result61[145]^and_result61[146]^and_result61[147]^and_result61[148]^and_result61[149]^and_result61[150]^and_result61[151]^and_result61[152]^and_result61[153]^and_result61[154]^and_result61[155]^and_result61[156]^and_result61[157]^and_result61[158]^and_result61[159]^and_result61[160]^and_result61[161]^and_result61[162]^and_result61[163]^and_result61[164]^and_result61[165]^and_result61[166]^and_result61[167]^and_result61[168]^and_result61[169]^and_result61[170]^and_result61[171]^and_result61[172]^and_result61[173]^and_result61[174]^and_result61[175]^and_result61[176]^and_result61[177]^and_result61[178]^and_result61[179]^and_result61[180]^and_result61[181]^and_result61[182]^and_result61[183]^and_result61[184]^and_result61[185]^and_result61[186]^and_result61[187]^and_result61[188]^and_result61[189]^and_result61[190]^and_result61[191]^and_result61[192]^and_result61[193]^and_result61[194]^and_result61[195]^and_result61[196]^and_result61[197]^and_result61[198]^and_result61[199]^and_result61[200]^and_result61[201]^and_result61[202]^and_result61[203]^and_result61[204]^and_result61[205]^and_result61[206]^and_result61[207]^and_result61[208]^and_result61[209]^and_result61[210]^and_result61[211]^and_result61[212]^and_result61[213]^and_result61[214]^and_result61[215]^and_result61[216]^and_result61[217]^and_result61[218]^and_result61[219]^and_result61[220]^and_result61[221]^and_result61[222]^and_result61[223]^and_result61[224]^and_result61[225]^and_result61[226]^and_result61[227]^and_result61[228]^and_result61[229]^and_result61[230]^and_result61[231]^and_result61[232]^and_result61[233]^and_result61[234]^and_result61[235]^and_result61[236]^and_result61[237]^and_result61[238]^and_result61[239]^and_result61[240]^and_result61[241]^and_result61[242]^and_result61[243]^and_result61[244]^and_result61[245]^and_result61[246]^and_result61[247]^and_result61[248]^and_result61[249]^and_result61[250]^and_result61[251]^and_result61[252]^and_result61[253]^and_result61[254];
assign key[62]=and_result62[0]^and_result62[1]^and_result62[2]^and_result62[3]^and_result62[4]^and_result62[5]^and_result62[6]^and_result62[7]^and_result62[8]^and_result62[9]^and_result62[10]^and_result62[11]^and_result62[12]^and_result62[13]^and_result62[14]^and_result62[15]^and_result62[16]^and_result62[17]^and_result62[18]^and_result62[19]^and_result62[20]^and_result62[21]^and_result62[22]^and_result62[23]^and_result62[24]^and_result62[25]^and_result62[26]^and_result62[27]^and_result62[28]^and_result62[29]^and_result62[30]^and_result62[31]^and_result62[32]^and_result62[33]^and_result62[34]^and_result62[35]^and_result62[36]^and_result62[37]^and_result62[38]^and_result62[39]^and_result62[40]^and_result62[41]^and_result62[42]^and_result62[43]^and_result62[44]^and_result62[45]^and_result62[46]^and_result62[47]^and_result62[48]^and_result62[49]^and_result62[50]^and_result62[51]^and_result62[52]^and_result62[53]^and_result62[54]^and_result62[55]^and_result62[56]^and_result62[57]^and_result62[58]^and_result62[59]^and_result62[60]^and_result62[61]^and_result62[62]^and_result62[63]^and_result62[64]^and_result62[65]^and_result62[66]^and_result62[67]^and_result62[68]^and_result62[69]^and_result62[70]^and_result62[71]^and_result62[72]^and_result62[73]^and_result62[74]^and_result62[75]^and_result62[76]^and_result62[77]^and_result62[78]^and_result62[79]^and_result62[80]^and_result62[81]^and_result62[82]^and_result62[83]^and_result62[84]^and_result62[85]^and_result62[86]^and_result62[87]^and_result62[88]^and_result62[89]^and_result62[90]^and_result62[91]^and_result62[92]^and_result62[93]^and_result62[94]^and_result62[95]^and_result62[96]^and_result62[97]^and_result62[98]^and_result62[99]^and_result62[100]^and_result62[101]^and_result62[102]^and_result62[103]^and_result62[104]^and_result62[105]^and_result62[106]^and_result62[107]^and_result62[108]^and_result62[109]^and_result62[110]^and_result62[111]^and_result62[112]^and_result62[113]^and_result62[114]^and_result62[115]^and_result62[116]^and_result62[117]^and_result62[118]^and_result62[119]^and_result62[120]^and_result62[121]^and_result62[122]^and_result62[123]^and_result62[124]^and_result62[125]^and_result62[126]^and_result62[127]^and_result62[128]^and_result62[129]^and_result62[130]^and_result62[131]^and_result62[132]^and_result62[133]^and_result62[134]^and_result62[135]^and_result62[136]^and_result62[137]^and_result62[138]^and_result62[139]^and_result62[140]^and_result62[141]^and_result62[142]^and_result62[143]^and_result62[144]^and_result62[145]^and_result62[146]^and_result62[147]^and_result62[148]^and_result62[149]^and_result62[150]^and_result62[151]^and_result62[152]^and_result62[153]^and_result62[154]^and_result62[155]^and_result62[156]^and_result62[157]^and_result62[158]^and_result62[159]^and_result62[160]^and_result62[161]^and_result62[162]^and_result62[163]^and_result62[164]^and_result62[165]^and_result62[166]^and_result62[167]^and_result62[168]^and_result62[169]^and_result62[170]^and_result62[171]^and_result62[172]^and_result62[173]^and_result62[174]^and_result62[175]^and_result62[176]^and_result62[177]^and_result62[178]^and_result62[179]^and_result62[180]^and_result62[181]^and_result62[182]^and_result62[183]^and_result62[184]^and_result62[185]^and_result62[186]^and_result62[187]^and_result62[188]^and_result62[189]^and_result62[190]^and_result62[191]^and_result62[192]^and_result62[193]^and_result62[194]^and_result62[195]^and_result62[196]^and_result62[197]^and_result62[198]^and_result62[199]^and_result62[200]^and_result62[201]^and_result62[202]^and_result62[203]^and_result62[204]^and_result62[205]^and_result62[206]^and_result62[207]^and_result62[208]^and_result62[209]^and_result62[210]^and_result62[211]^and_result62[212]^and_result62[213]^and_result62[214]^and_result62[215]^and_result62[216]^and_result62[217]^and_result62[218]^and_result62[219]^and_result62[220]^and_result62[221]^and_result62[222]^and_result62[223]^and_result62[224]^and_result62[225]^and_result62[226]^and_result62[227]^and_result62[228]^and_result62[229]^and_result62[230]^and_result62[231]^and_result62[232]^and_result62[233]^and_result62[234]^and_result62[235]^and_result62[236]^and_result62[237]^and_result62[238]^and_result62[239]^and_result62[240]^and_result62[241]^and_result62[242]^and_result62[243]^and_result62[244]^and_result62[245]^and_result62[246]^and_result62[247]^and_result62[248]^and_result62[249]^and_result62[250]^and_result62[251]^and_result62[252]^and_result62[253]^and_result62[254];
assign key[63]=and_result63[0]^and_result63[1]^and_result63[2]^and_result63[3]^and_result63[4]^and_result63[5]^and_result63[6]^and_result63[7]^and_result63[8]^and_result63[9]^and_result63[10]^and_result63[11]^and_result63[12]^and_result63[13]^and_result63[14]^and_result63[15]^and_result63[16]^and_result63[17]^and_result63[18]^and_result63[19]^and_result63[20]^and_result63[21]^and_result63[22]^and_result63[23]^and_result63[24]^and_result63[25]^and_result63[26]^and_result63[27]^and_result63[28]^and_result63[29]^and_result63[30]^and_result63[31]^and_result63[32]^and_result63[33]^and_result63[34]^and_result63[35]^and_result63[36]^and_result63[37]^and_result63[38]^and_result63[39]^and_result63[40]^and_result63[41]^and_result63[42]^and_result63[43]^and_result63[44]^and_result63[45]^and_result63[46]^and_result63[47]^and_result63[48]^and_result63[49]^and_result63[50]^and_result63[51]^and_result63[52]^and_result63[53]^and_result63[54]^and_result63[55]^and_result63[56]^and_result63[57]^and_result63[58]^and_result63[59]^and_result63[60]^and_result63[61]^and_result63[62]^and_result63[63]^and_result63[64]^and_result63[65]^and_result63[66]^and_result63[67]^and_result63[68]^and_result63[69]^and_result63[70]^and_result63[71]^and_result63[72]^and_result63[73]^and_result63[74]^and_result63[75]^and_result63[76]^and_result63[77]^and_result63[78]^and_result63[79]^and_result63[80]^and_result63[81]^and_result63[82]^and_result63[83]^and_result63[84]^and_result63[85]^and_result63[86]^and_result63[87]^and_result63[88]^and_result63[89]^and_result63[90]^and_result63[91]^and_result63[92]^and_result63[93]^and_result63[94]^and_result63[95]^and_result63[96]^and_result63[97]^and_result63[98]^and_result63[99]^and_result63[100]^and_result63[101]^and_result63[102]^and_result63[103]^and_result63[104]^and_result63[105]^and_result63[106]^and_result63[107]^and_result63[108]^and_result63[109]^and_result63[110]^and_result63[111]^and_result63[112]^and_result63[113]^and_result63[114]^and_result63[115]^and_result63[116]^and_result63[117]^and_result63[118]^and_result63[119]^and_result63[120]^and_result63[121]^and_result63[122]^and_result63[123]^and_result63[124]^and_result63[125]^and_result63[126]^and_result63[127]^and_result63[128]^and_result63[129]^and_result63[130]^and_result63[131]^and_result63[132]^and_result63[133]^and_result63[134]^and_result63[135]^and_result63[136]^and_result63[137]^and_result63[138]^and_result63[139]^and_result63[140]^and_result63[141]^and_result63[142]^and_result63[143]^and_result63[144]^and_result63[145]^and_result63[146]^and_result63[147]^and_result63[148]^and_result63[149]^and_result63[150]^and_result63[151]^and_result63[152]^and_result63[153]^and_result63[154]^and_result63[155]^and_result63[156]^and_result63[157]^and_result63[158]^and_result63[159]^and_result63[160]^and_result63[161]^and_result63[162]^and_result63[163]^and_result63[164]^and_result63[165]^and_result63[166]^and_result63[167]^and_result63[168]^and_result63[169]^and_result63[170]^and_result63[171]^and_result63[172]^and_result63[173]^and_result63[174]^and_result63[175]^and_result63[176]^and_result63[177]^and_result63[178]^and_result63[179]^and_result63[180]^and_result63[181]^and_result63[182]^and_result63[183]^and_result63[184]^and_result63[185]^and_result63[186]^and_result63[187]^and_result63[188]^and_result63[189]^and_result63[190]^and_result63[191]^and_result63[192]^and_result63[193]^and_result63[194]^and_result63[195]^and_result63[196]^and_result63[197]^and_result63[198]^and_result63[199]^and_result63[200]^and_result63[201]^and_result63[202]^and_result63[203]^and_result63[204]^and_result63[205]^and_result63[206]^and_result63[207]^and_result63[208]^and_result63[209]^and_result63[210]^and_result63[211]^and_result63[212]^and_result63[213]^and_result63[214]^and_result63[215]^and_result63[216]^and_result63[217]^and_result63[218]^and_result63[219]^and_result63[220]^and_result63[221]^and_result63[222]^and_result63[223]^and_result63[224]^and_result63[225]^and_result63[226]^and_result63[227]^and_result63[228]^and_result63[229]^and_result63[230]^and_result63[231]^and_result63[232]^and_result63[233]^and_result63[234]^and_result63[235]^and_result63[236]^and_result63[237]^and_result63[238]^and_result63[239]^and_result63[240]^and_result63[241]^and_result63[242]^and_result63[243]^and_result63[244]^and_result63[245]^and_result63[246]^and_result63[247]^and_result63[248]^and_result63[249]^and_result63[250]^and_result63[251]^and_result63[252]^and_result63[253]^and_result63[254];
assign key[64]=and_result64[0]^and_result64[1]^and_result64[2]^and_result64[3]^and_result64[4]^and_result64[5]^and_result64[6]^and_result64[7]^and_result64[8]^and_result64[9]^and_result64[10]^and_result64[11]^and_result64[12]^and_result64[13]^and_result64[14]^and_result64[15]^and_result64[16]^and_result64[17]^and_result64[18]^and_result64[19]^and_result64[20]^and_result64[21]^and_result64[22]^and_result64[23]^and_result64[24]^and_result64[25]^and_result64[26]^and_result64[27]^and_result64[28]^and_result64[29]^and_result64[30]^and_result64[31]^and_result64[32]^and_result64[33]^and_result64[34]^and_result64[35]^and_result64[36]^and_result64[37]^and_result64[38]^and_result64[39]^and_result64[40]^and_result64[41]^and_result64[42]^and_result64[43]^and_result64[44]^and_result64[45]^and_result64[46]^and_result64[47]^and_result64[48]^and_result64[49]^and_result64[50]^and_result64[51]^and_result64[52]^and_result64[53]^and_result64[54]^and_result64[55]^and_result64[56]^and_result64[57]^and_result64[58]^and_result64[59]^and_result64[60]^and_result64[61]^and_result64[62]^and_result64[63]^and_result64[64]^and_result64[65]^and_result64[66]^and_result64[67]^and_result64[68]^and_result64[69]^and_result64[70]^and_result64[71]^and_result64[72]^and_result64[73]^and_result64[74]^and_result64[75]^and_result64[76]^and_result64[77]^and_result64[78]^and_result64[79]^and_result64[80]^and_result64[81]^and_result64[82]^and_result64[83]^and_result64[84]^and_result64[85]^and_result64[86]^and_result64[87]^and_result64[88]^and_result64[89]^and_result64[90]^and_result64[91]^and_result64[92]^and_result64[93]^and_result64[94]^and_result64[95]^and_result64[96]^and_result64[97]^and_result64[98]^and_result64[99]^and_result64[100]^and_result64[101]^and_result64[102]^and_result64[103]^and_result64[104]^and_result64[105]^and_result64[106]^and_result64[107]^and_result64[108]^and_result64[109]^and_result64[110]^and_result64[111]^and_result64[112]^and_result64[113]^and_result64[114]^and_result64[115]^and_result64[116]^and_result64[117]^and_result64[118]^and_result64[119]^and_result64[120]^and_result64[121]^and_result64[122]^and_result64[123]^and_result64[124]^and_result64[125]^and_result64[126]^and_result64[127]^and_result64[128]^and_result64[129]^and_result64[130]^and_result64[131]^and_result64[132]^and_result64[133]^and_result64[134]^and_result64[135]^and_result64[136]^and_result64[137]^and_result64[138]^and_result64[139]^and_result64[140]^and_result64[141]^and_result64[142]^and_result64[143]^and_result64[144]^and_result64[145]^and_result64[146]^and_result64[147]^and_result64[148]^and_result64[149]^and_result64[150]^and_result64[151]^and_result64[152]^and_result64[153]^and_result64[154]^and_result64[155]^and_result64[156]^and_result64[157]^and_result64[158]^and_result64[159]^and_result64[160]^and_result64[161]^and_result64[162]^and_result64[163]^and_result64[164]^and_result64[165]^and_result64[166]^and_result64[167]^and_result64[168]^and_result64[169]^and_result64[170]^and_result64[171]^and_result64[172]^and_result64[173]^and_result64[174]^and_result64[175]^and_result64[176]^and_result64[177]^and_result64[178]^and_result64[179]^and_result64[180]^and_result64[181]^and_result64[182]^and_result64[183]^and_result64[184]^and_result64[185]^and_result64[186]^and_result64[187]^and_result64[188]^and_result64[189]^and_result64[190]^and_result64[191]^and_result64[192]^and_result64[193]^and_result64[194]^and_result64[195]^and_result64[196]^and_result64[197]^and_result64[198]^and_result64[199]^and_result64[200]^and_result64[201]^and_result64[202]^and_result64[203]^and_result64[204]^and_result64[205]^and_result64[206]^and_result64[207]^and_result64[208]^and_result64[209]^and_result64[210]^and_result64[211]^and_result64[212]^and_result64[213]^and_result64[214]^and_result64[215]^and_result64[216]^and_result64[217]^and_result64[218]^and_result64[219]^and_result64[220]^and_result64[221]^and_result64[222]^and_result64[223]^and_result64[224]^and_result64[225]^and_result64[226]^and_result64[227]^and_result64[228]^and_result64[229]^and_result64[230]^and_result64[231]^and_result64[232]^and_result64[233]^and_result64[234]^and_result64[235]^and_result64[236]^and_result64[237]^and_result64[238]^and_result64[239]^and_result64[240]^and_result64[241]^and_result64[242]^and_result64[243]^and_result64[244]^and_result64[245]^and_result64[246]^and_result64[247]^and_result64[248]^and_result64[249]^and_result64[250]^and_result64[251]^and_result64[252]^and_result64[253]^and_result64[254];
assign key[65]=and_result65[0]^and_result65[1]^and_result65[2]^and_result65[3]^and_result65[4]^and_result65[5]^and_result65[6]^and_result65[7]^and_result65[8]^and_result65[9]^and_result65[10]^and_result65[11]^and_result65[12]^and_result65[13]^and_result65[14]^and_result65[15]^and_result65[16]^and_result65[17]^and_result65[18]^and_result65[19]^and_result65[20]^and_result65[21]^and_result65[22]^and_result65[23]^and_result65[24]^and_result65[25]^and_result65[26]^and_result65[27]^and_result65[28]^and_result65[29]^and_result65[30]^and_result65[31]^and_result65[32]^and_result65[33]^and_result65[34]^and_result65[35]^and_result65[36]^and_result65[37]^and_result65[38]^and_result65[39]^and_result65[40]^and_result65[41]^and_result65[42]^and_result65[43]^and_result65[44]^and_result65[45]^and_result65[46]^and_result65[47]^and_result65[48]^and_result65[49]^and_result65[50]^and_result65[51]^and_result65[52]^and_result65[53]^and_result65[54]^and_result65[55]^and_result65[56]^and_result65[57]^and_result65[58]^and_result65[59]^and_result65[60]^and_result65[61]^and_result65[62]^and_result65[63]^and_result65[64]^and_result65[65]^and_result65[66]^and_result65[67]^and_result65[68]^and_result65[69]^and_result65[70]^and_result65[71]^and_result65[72]^and_result65[73]^and_result65[74]^and_result65[75]^and_result65[76]^and_result65[77]^and_result65[78]^and_result65[79]^and_result65[80]^and_result65[81]^and_result65[82]^and_result65[83]^and_result65[84]^and_result65[85]^and_result65[86]^and_result65[87]^and_result65[88]^and_result65[89]^and_result65[90]^and_result65[91]^and_result65[92]^and_result65[93]^and_result65[94]^and_result65[95]^and_result65[96]^and_result65[97]^and_result65[98]^and_result65[99]^and_result65[100]^and_result65[101]^and_result65[102]^and_result65[103]^and_result65[104]^and_result65[105]^and_result65[106]^and_result65[107]^and_result65[108]^and_result65[109]^and_result65[110]^and_result65[111]^and_result65[112]^and_result65[113]^and_result65[114]^and_result65[115]^and_result65[116]^and_result65[117]^and_result65[118]^and_result65[119]^and_result65[120]^and_result65[121]^and_result65[122]^and_result65[123]^and_result65[124]^and_result65[125]^and_result65[126]^and_result65[127]^and_result65[128]^and_result65[129]^and_result65[130]^and_result65[131]^and_result65[132]^and_result65[133]^and_result65[134]^and_result65[135]^and_result65[136]^and_result65[137]^and_result65[138]^and_result65[139]^and_result65[140]^and_result65[141]^and_result65[142]^and_result65[143]^and_result65[144]^and_result65[145]^and_result65[146]^and_result65[147]^and_result65[148]^and_result65[149]^and_result65[150]^and_result65[151]^and_result65[152]^and_result65[153]^and_result65[154]^and_result65[155]^and_result65[156]^and_result65[157]^and_result65[158]^and_result65[159]^and_result65[160]^and_result65[161]^and_result65[162]^and_result65[163]^and_result65[164]^and_result65[165]^and_result65[166]^and_result65[167]^and_result65[168]^and_result65[169]^and_result65[170]^and_result65[171]^and_result65[172]^and_result65[173]^and_result65[174]^and_result65[175]^and_result65[176]^and_result65[177]^and_result65[178]^and_result65[179]^and_result65[180]^and_result65[181]^and_result65[182]^and_result65[183]^and_result65[184]^and_result65[185]^and_result65[186]^and_result65[187]^and_result65[188]^and_result65[189]^and_result65[190]^and_result65[191]^and_result65[192]^and_result65[193]^and_result65[194]^and_result65[195]^and_result65[196]^and_result65[197]^and_result65[198]^and_result65[199]^and_result65[200]^and_result65[201]^and_result65[202]^and_result65[203]^and_result65[204]^and_result65[205]^and_result65[206]^and_result65[207]^and_result65[208]^and_result65[209]^and_result65[210]^and_result65[211]^and_result65[212]^and_result65[213]^and_result65[214]^and_result65[215]^and_result65[216]^and_result65[217]^and_result65[218]^and_result65[219]^and_result65[220]^and_result65[221]^and_result65[222]^and_result65[223]^and_result65[224]^and_result65[225]^and_result65[226]^and_result65[227]^and_result65[228]^and_result65[229]^and_result65[230]^and_result65[231]^and_result65[232]^and_result65[233]^and_result65[234]^and_result65[235]^and_result65[236]^and_result65[237]^and_result65[238]^and_result65[239]^and_result65[240]^and_result65[241]^and_result65[242]^and_result65[243]^and_result65[244]^and_result65[245]^and_result65[246]^and_result65[247]^and_result65[248]^and_result65[249]^and_result65[250]^and_result65[251]^and_result65[252]^and_result65[253]^and_result65[254];
assign key[66]=and_result66[0]^and_result66[1]^and_result66[2]^and_result66[3]^and_result66[4]^and_result66[5]^and_result66[6]^and_result66[7]^and_result66[8]^and_result66[9]^and_result66[10]^and_result66[11]^and_result66[12]^and_result66[13]^and_result66[14]^and_result66[15]^and_result66[16]^and_result66[17]^and_result66[18]^and_result66[19]^and_result66[20]^and_result66[21]^and_result66[22]^and_result66[23]^and_result66[24]^and_result66[25]^and_result66[26]^and_result66[27]^and_result66[28]^and_result66[29]^and_result66[30]^and_result66[31]^and_result66[32]^and_result66[33]^and_result66[34]^and_result66[35]^and_result66[36]^and_result66[37]^and_result66[38]^and_result66[39]^and_result66[40]^and_result66[41]^and_result66[42]^and_result66[43]^and_result66[44]^and_result66[45]^and_result66[46]^and_result66[47]^and_result66[48]^and_result66[49]^and_result66[50]^and_result66[51]^and_result66[52]^and_result66[53]^and_result66[54]^and_result66[55]^and_result66[56]^and_result66[57]^and_result66[58]^and_result66[59]^and_result66[60]^and_result66[61]^and_result66[62]^and_result66[63]^and_result66[64]^and_result66[65]^and_result66[66]^and_result66[67]^and_result66[68]^and_result66[69]^and_result66[70]^and_result66[71]^and_result66[72]^and_result66[73]^and_result66[74]^and_result66[75]^and_result66[76]^and_result66[77]^and_result66[78]^and_result66[79]^and_result66[80]^and_result66[81]^and_result66[82]^and_result66[83]^and_result66[84]^and_result66[85]^and_result66[86]^and_result66[87]^and_result66[88]^and_result66[89]^and_result66[90]^and_result66[91]^and_result66[92]^and_result66[93]^and_result66[94]^and_result66[95]^and_result66[96]^and_result66[97]^and_result66[98]^and_result66[99]^and_result66[100]^and_result66[101]^and_result66[102]^and_result66[103]^and_result66[104]^and_result66[105]^and_result66[106]^and_result66[107]^and_result66[108]^and_result66[109]^and_result66[110]^and_result66[111]^and_result66[112]^and_result66[113]^and_result66[114]^and_result66[115]^and_result66[116]^and_result66[117]^and_result66[118]^and_result66[119]^and_result66[120]^and_result66[121]^and_result66[122]^and_result66[123]^and_result66[124]^and_result66[125]^and_result66[126]^and_result66[127]^and_result66[128]^and_result66[129]^and_result66[130]^and_result66[131]^and_result66[132]^and_result66[133]^and_result66[134]^and_result66[135]^and_result66[136]^and_result66[137]^and_result66[138]^and_result66[139]^and_result66[140]^and_result66[141]^and_result66[142]^and_result66[143]^and_result66[144]^and_result66[145]^and_result66[146]^and_result66[147]^and_result66[148]^and_result66[149]^and_result66[150]^and_result66[151]^and_result66[152]^and_result66[153]^and_result66[154]^and_result66[155]^and_result66[156]^and_result66[157]^and_result66[158]^and_result66[159]^and_result66[160]^and_result66[161]^and_result66[162]^and_result66[163]^and_result66[164]^and_result66[165]^and_result66[166]^and_result66[167]^and_result66[168]^and_result66[169]^and_result66[170]^and_result66[171]^and_result66[172]^and_result66[173]^and_result66[174]^and_result66[175]^and_result66[176]^and_result66[177]^and_result66[178]^and_result66[179]^and_result66[180]^and_result66[181]^and_result66[182]^and_result66[183]^and_result66[184]^and_result66[185]^and_result66[186]^and_result66[187]^and_result66[188]^and_result66[189]^and_result66[190]^and_result66[191]^and_result66[192]^and_result66[193]^and_result66[194]^and_result66[195]^and_result66[196]^and_result66[197]^and_result66[198]^and_result66[199]^and_result66[200]^and_result66[201]^and_result66[202]^and_result66[203]^and_result66[204]^and_result66[205]^and_result66[206]^and_result66[207]^and_result66[208]^and_result66[209]^and_result66[210]^and_result66[211]^and_result66[212]^and_result66[213]^and_result66[214]^and_result66[215]^and_result66[216]^and_result66[217]^and_result66[218]^and_result66[219]^and_result66[220]^and_result66[221]^and_result66[222]^and_result66[223]^and_result66[224]^and_result66[225]^and_result66[226]^and_result66[227]^and_result66[228]^and_result66[229]^and_result66[230]^and_result66[231]^and_result66[232]^and_result66[233]^and_result66[234]^and_result66[235]^and_result66[236]^and_result66[237]^and_result66[238]^and_result66[239]^and_result66[240]^and_result66[241]^and_result66[242]^and_result66[243]^and_result66[244]^and_result66[245]^and_result66[246]^and_result66[247]^and_result66[248]^and_result66[249]^and_result66[250]^and_result66[251]^and_result66[252]^and_result66[253]^and_result66[254];
assign key[67]=and_result67[0]^and_result67[1]^and_result67[2]^and_result67[3]^and_result67[4]^and_result67[5]^and_result67[6]^and_result67[7]^and_result67[8]^and_result67[9]^and_result67[10]^and_result67[11]^and_result67[12]^and_result67[13]^and_result67[14]^and_result67[15]^and_result67[16]^and_result67[17]^and_result67[18]^and_result67[19]^and_result67[20]^and_result67[21]^and_result67[22]^and_result67[23]^and_result67[24]^and_result67[25]^and_result67[26]^and_result67[27]^and_result67[28]^and_result67[29]^and_result67[30]^and_result67[31]^and_result67[32]^and_result67[33]^and_result67[34]^and_result67[35]^and_result67[36]^and_result67[37]^and_result67[38]^and_result67[39]^and_result67[40]^and_result67[41]^and_result67[42]^and_result67[43]^and_result67[44]^and_result67[45]^and_result67[46]^and_result67[47]^and_result67[48]^and_result67[49]^and_result67[50]^and_result67[51]^and_result67[52]^and_result67[53]^and_result67[54]^and_result67[55]^and_result67[56]^and_result67[57]^and_result67[58]^and_result67[59]^and_result67[60]^and_result67[61]^and_result67[62]^and_result67[63]^and_result67[64]^and_result67[65]^and_result67[66]^and_result67[67]^and_result67[68]^and_result67[69]^and_result67[70]^and_result67[71]^and_result67[72]^and_result67[73]^and_result67[74]^and_result67[75]^and_result67[76]^and_result67[77]^and_result67[78]^and_result67[79]^and_result67[80]^and_result67[81]^and_result67[82]^and_result67[83]^and_result67[84]^and_result67[85]^and_result67[86]^and_result67[87]^and_result67[88]^and_result67[89]^and_result67[90]^and_result67[91]^and_result67[92]^and_result67[93]^and_result67[94]^and_result67[95]^and_result67[96]^and_result67[97]^and_result67[98]^and_result67[99]^and_result67[100]^and_result67[101]^and_result67[102]^and_result67[103]^and_result67[104]^and_result67[105]^and_result67[106]^and_result67[107]^and_result67[108]^and_result67[109]^and_result67[110]^and_result67[111]^and_result67[112]^and_result67[113]^and_result67[114]^and_result67[115]^and_result67[116]^and_result67[117]^and_result67[118]^and_result67[119]^and_result67[120]^and_result67[121]^and_result67[122]^and_result67[123]^and_result67[124]^and_result67[125]^and_result67[126]^and_result67[127]^and_result67[128]^and_result67[129]^and_result67[130]^and_result67[131]^and_result67[132]^and_result67[133]^and_result67[134]^and_result67[135]^and_result67[136]^and_result67[137]^and_result67[138]^and_result67[139]^and_result67[140]^and_result67[141]^and_result67[142]^and_result67[143]^and_result67[144]^and_result67[145]^and_result67[146]^and_result67[147]^and_result67[148]^and_result67[149]^and_result67[150]^and_result67[151]^and_result67[152]^and_result67[153]^and_result67[154]^and_result67[155]^and_result67[156]^and_result67[157]^and_result67[158]^and_result67[159]^and_result67[160]^and_result67[161]^and_result67[162]^and_result67[163]^and_result67[164]^and_result67[165]^and_result67[166]^and_result67[167]^and_result67[168]^and_result67[169]^and_result67[170]^and_result67[171]^and_result67[172]^and_result67[173]^and_result67[174]^and_result67[175]^and_result67[176]^and_result67[177]^and_result67[178]^and_result67[179]^and_result67[180]^and_result67[181]^and_result67[182]^and_result67[183]^and_result67[184]^and_result67[185]^and_result67[186]^and_result67[187]^and_result67[188]^and_result67[189]^and_result67[190]^and_result67[191]^and_result67[192]^and_result67[193]^and_result67[194]^and_result67[195]^and_result67[196]^and_result67[197]^and_result67[198]^and_result67[199]^and_result67[200]^and_result67[201]^and_result67[202]^and_result67[203]^and_result67[204]^and_result67[205]^and_result67[206]^and_result67[207]^and_result67[208]^and_result67[209]^and_result67[210]^and_result67[211]^and_result67[212]^and_result67[213]^and_result67[214]^and_result67[215]^and_result67[216]^and_result67[217]^and_result67[218]^and_result67[219]^and_result67[220]^and_result67[221]^and_result67[222]^and_result67[223]^and_result67[224]^and_result67[225]^and_result67[226]^and_result67[227]^and_result67[228]^and_result67[229]^and_result67[230]^and_result67[231]^and_result67[232]^and_result67[233]^and_result67[234]^and_result67[235]^and_result67[236]^and_result67[237]^and_result67[238]^and_result67[239]^and_result67[240]^and_result67[241]^and_result67[242]^and_result67[243]^and_result67[244]^and_result67[245]^and_result67[246]^and_result67[247]^and_result67[248]^and_result67[249]^and_result67[250]^and_result67[251]^and_result67[252]^and_result67[253]^and_result67[254];
assign key[68]=and_result68[0]^and_result68[1]^and_result68[2]^and_result68[3]^and_result68[4]^and_result68[5]^and_result68[6]^and_result68[7]^and_result68[8]^and_result68[9]^and_result68[10]^and_result68[11]^and_result68[12]^and_result68[13]^and_result68[14]^and_result68[15]^and_result68[16]^and_result68[17]^and_result68[18]^and_result68[19]^and_result68[20]^and_result68[21]^and_result68[22]^and_result68[23]^and_result68[24]^and_result68[25]^and_result68[26]^and_result68[27]^and_result68[28]^and_result68[29]^and_result68[30]^and_result68[31]^and_result68[32]^and_result68[33]^and_result68[34]^and_result68[35]^and_result68[36]^and_result68[37]^and_result68[38]^and_result68[39]^and_result68[40]^and_result68[41]^and_result68[42]^and_result68[43]^and_result68[44]^and_result68[45]^and_result68[46]^and_result68[47]^and_result68[48]^and_result68[49]^and_result68[50]^and_result68[51]^and_result68[52]^and_result68[53]^and_result68[54]^and_result68[55]^and_result68[56]^and_result68[57]^and_result68[58]^and_result68[59]^and_result68[60]^and_result68[61]^and_result68[62]^and_result68[63]^and_result68[64]^and_result68[65]^and_result68[66]^and_result68[67]^and_result68[68]^and_result68[69]^and_result68[70]^and_result68[71]^and_result68[72]^and_result68[73]^and_result68[74]^and_result68[75]^and_result68[76]^and_result68[77]^and_result68[78]^and_result68[79]^and_result68[80]^and_result68[81]^and_result68[82]^and_result68[83]^and_result68[84]^and_result68[85]^and_result68[86]^and_result68[87]^and_result68[88]^and_result68[89]^and_result68[90]^and_result68[91]^and_result68[92]^and_result68[93]^and_result68[94]^and_result68[95]^and_result68[96]^and_result68[97]^and_result68[98]^and_result68[99]^and_result68[100]^and_result68[101]^and_result68[102]^and_result68[103]^and_result68[104]^and_result68[105]^and_result68[106]^and_result68[107]^and_result68[108]^and_result68[109]^and_result68[110]^and_result68[111]^and_result68[112]^and_result68[113]^and_result68[114]^and_result68[115]^and_result68[116]^and_result68[117]^and_result68[118]^and_result68[119]^and_result68[120]^and_result68[121]^and_result68[122]^and_result68[123]^and_result68[124]^and_result68[125]^and_result68[126]^and_result68[127]^and_result68[128]^and_result68[129]^and_result68[130]^and_result68[131]^and_result68[132]^and_result68[133]^and_result68[134]^and_result68[135]^and_result68[136]^and_result68[137]^and_result68[138]^and_result68[139]^and_result68[140]^and_result68[141]^and_result68[142]^and_result68[143]^and_result68[144]^and_result68[145]^and_result68[146]^and_result68[147]^and_result68[148]^and_result68[149]^and_result68[150]^and_result68[151]^and_result68[152]^and_result68[153]^and_result68[154]^and_result68[155]^and_result68[156]^and_result68[157]^and_result68[158]^and_result68[159]^and_result68[160]^and_result68[161]^and_result68[162]^and_result68[163]^and_result68[164]^and_result68[165]^and_result68[166]^and_result68[167]^and_result68[168]^and_result68[169]^and_result68[170]^and_result68[171]^and_result68[172]^and_result68[173]^and_result68[174]^and_result68[175]^and_result68[176]^and_result68[177]^and_result68[178]^and_result68[179]^and_result68[180]^and_result68[181]^and_result68[182]^and_result68[183]^and_result68[184]^and_result68[185]^and_result68[186]^and_result68[187]^and_result68[188]^and_result68[189]^and_result68[190]^and_result68[191]^and_result68[192]^and_result68[193]^and_result68[194]^and_result68[195]^and_result68[196]^and_result68[197]^and_result68[198]^and_result68[199]^and_result68[200]^and_result68[201]^and_result68[202]^and_result68[203]^and_result68[204]^and_result68[205]^and_result68[206]^and_result68[207]^and_result68[208]^and_result68[209]^and_result68[210]^and_result68[211]^and_result68[212]^and_result68[213]^and_result68[214]^and_result68[215]^and_result68[216]^and_result68[217]^and_result68[218]^and_result68[219]^and_result68[220]^and_result68[221]^and_result68[222]^and_result68[223]^and_result68[224]^and_result68[225]^and_result68[226]^and_result68[227]^and_result68[228]^and_result68[229]^and_result68[230]^and_result68[231]^and_result68[232]^and_result68[233]^and_result68[234]^and_result68[235]^and_result68[236]^and_result68[237]^and_result68[238]^and_result68[239]^and_result68[240]^and_result68[241]^and_result68[242]^and_result68[243]^and_result68[244]^and_result68[245]^and_result68[246]^and_result68[247]^and_result68[248]^and_result68[249]^and_result68[250]^and_result68[251]^and_result68[252]^and_result68[253]^and_result68[254];
assign key[69]=and_result69[0]^and_result69[1]^and_result69[2]^and_result69[3]^and_result69[4]^and_result69[5]^and_result69[6]^and_result69[7]^and_result69[8]^and_result69[9]^and_result69[10]^and_result69[11]^and_result69[12]^and_result69[13]^and_result69[14]^and_result69[15]^and_result69[16]^and_result69[17]^and_result69[18]^and_result69[19]^and_result69[20]^and_result69[21]^and_result69[22]^and_result69[23]^and_result69[24]^and_result69[25]^and_result69[26]^and_result69[27]^and_result69[28]^and_result69[29]^and_result69[30]^and_result69[31]^and_result69[32]^and_result69[33]^and_result69[34]^and_result69[35]^and_result69[36]^and_result69[37]^and_result69[38]^and_result69[39]^and_result69[40]^and_result69[41]^and_result69[42]^and_result69[43]^and_result69[44]^and_result69[45]^and_result69[46]^and_result69[47]^and_result69[48]^and_result69[49]^and_result69[50]^and_result69[51]^and_result69[52]^and_result69[53]^and_result69[54]^and_result69[55]^and_result69[56]^and_result69[57]^and_result69[58]^and_result69[59]^and_result69[60]^and_result69[61]^and_result69[62]^and_result69[63]^and_result69[64]^and_result69[65]^and_result69[66]^and_result69[67]^and_result69[68]^and_result69[69]^and_result69[70]^and_result69[71]^and_result69[72]^and_result69[73]^and_result69[74]^and_result69[75]^and_result69[76]^and_result69[77]^and_result69[78]^and_result69[79]^and_result69[80]^and_result69[81]^and_result69[82]^and_result69[83]^and_result69[84]^and_result69[85]^and_result69[86]^and_result69[87]^and_result69[88]^and_result69[89]^and_result69[90]^and_result69[91]^and_result69[92]^and_result69[93]^and_result69[94]^and_result69[95]^and_result69[96]^and_result69[97]^and_result69[98]^and_result69[99]^and_result69[100]^and_result69[101]^and_result69[102]^and_result69[103]^and_result69[104]^and_result69[105]^and_result69[106]^and_result69[107]^and_result69[108]^and_result69[109]^and_result69[110]^and_result69[111]^and_result69[112]^and_result69[113]^and_result69[114]^and_result69[115]^and_result69[116]^and_result69[117]^and_result69[118]^and_result69[119]^and_result69[120]^and_result69[121]^and_result69[122]^and_result69[123]^and_result69[124]^and_result69[125]^and_result69[126]^and_result69[127]^and_result69[128]^and_result69[129]^and_result69[130]^and_result69[131]^and_result69[132]^and_result69[133]^and_result69[134]^and_result69[135]^and_result69[136]^and_result69[137]^and_result69[138]^and_result69[139]^and_result69[140]^and_result69[141]^and_result69[142]^and_result69[143]^and_result69[144]^and_result69[145]^and_result69[146]^and_result69[147]^and_result69[148]^and_result69[149]^and_result69[150]^and_result69[151]^and_result69[152]^and_result69[153]^and_result69[154]^and_result69[155]^and_result69[156]^and_result69[157]^and_result69[158]^and_result69[159]^and_result69[160]^and_result69[161]^and_result69[162]^and_result69[163]^and_result69[164]^and_result69[165]^and_result69[166]^and_result69[167]^and_result69[168]^and_result69[169]^and_result69[170]^and_result69[171]^and_result69[172]^and_result69[173]^and_result69[174]^and_result69[175]^and_result69[176]^and_result69[177]^and_result69[178]^and_result69[179]^and_result69[180]^and_result69[181]^and_result69[182]^and_result69[183]^and_result69[184]^and_result69[185]^and_result69[186]^and_result69[187]^and_result69[188]^and_result69[189]^and_result69[190]^and_result69[191]^and_result69[192]^and_result69[193]^and_result69[194]^and_result69[195]^and_result69[196]^and_result69[197]^and_result69[198]^and_result69[199]^and_result69[200]^and_result69[201]^and_result69[202]^and_result69[203]^and_result69[204]^and_result69[205]^and_result69[206]^and_result69[207]^and_result69[208]^and_result69[209]^and_result69[210]^and_result69[211]^and_result69[212]^and_result69[213]^and_result69[214]^and_result69[215]^and_result69[216]^and_result69[217]^and_result69[218]^and_result69[219]^and_result69[220]^and_result69[221]^and_result69[222]^and_result69[223]^and_result69[224]^and_result69[225]^and_result69[226]^and_result69[227]^and_result69[228]^and_result69[229]^and_result69[230]^and_result69[231]^and_result69[232]^and_result69[233]^and_result69[234]^and_result69[235]^and_result69[236]^and_result69[237]^and_result69[238]^and_result69[239]^and_result69[240]^and_result69[241]^and_result69[242]^and_result69[243]^and_result69[244]^and_result69[245]^and_result69[246]^and_result69[247]^and_result69[248]^and_result69[249]^and_result69[250]^and_result69[251]^and_result69[252]^and_result69[253]^and_result69[254];
assign key[70]=and_result70[0]^and_result70[1]^and_result70[2]^and_result70[3]^and_result70[4]^and_result70[5]^and_result70[6]^and_result70[7]^and_result70[8]^and_result70[9]^and_result70[10]^and_result70[11]^and_result70[12]^and_result70[13]^and_result70[14]^and_result70[15]^and_result70[16]^and_result70[17]^and_result70[18]^and_result70[19]^and_result70[20]^and_result70[21]^and_result70[22]^and_result70[23]^and_result70[24]^and_result70[25]^and_result70[26]^and_result70[27]^and_result70[28]^and_result70[29]^and_result70[30]^and_result70[31]^and_result70[32]^and_result70[33]^and_result70[34]^and_result70[35]^and_result70[36]^and_result70[37]^and_result70[38]^and_result70[39]^and_result70[40]^and_result70[41]^and_result70[42]^and_result70[43]^and_result70[44]^and_result70[45]^and_result70[46]^and_result70[47]^and_result70[48]^and_result70[49]^and_result70[50]^and_result70[51]^and_result70[52]^and_result70[53]^and_result70[54]^and_result70[55]^and_result70[56]^and_result70[57]^and_result70[58]^and_result70[59]^and_result70[60]^and_result70[61]^and_result70[62]^and_result70[63]^and_result70[64]^and_result70[65]^and_result70[66]^and_result70[67]^and_result70[68]^and_result70[69]^and_result70[70]^and_result70[71]^and_result70[72]^and_result70[73]^and_result70[74]^and_result70[75]^and_result70[76]^and_result70[77]^and_result70[78]^and_result70[79]^and_result70[80]^and_result70[81]^and_result70[82]^and_result70[83]^and_result70[84]^and_result70[85]^and_result70[86]^and_result70[87]^and_result70[88]^and_result70[89]^and_result70[90]^and_result70[91]^and_result70[92]^and_result70[93]^and_result70[94]^and_result70[95]^and_result70[96]^and_result70[97]^and_result70[98]^and_result70[99]^and_result70[100]^and_result70[101]^and_result70[102]^and_result70[103]^and_result70[104]^and_result70[105]^and_result70[106]^and_result70[107]^and_result70[108]^and_result70[109]^and_result70[110]^and_result70[111]^and_result70[112]^and_result70[113]^and_result70[114]^and_result70[115]^and_result70[116]^and_result70[117]^and_result70[118]^and_result70[119]^and_result70[120]^and_result70[121]^and_result70[122]^and_result70[123]^and_result70[124]^and_result70[125]^and_result70[126]^and_result70[127]^and_result70[128]^and_result70[129]^and_result70[130]^and_result70[131]^and_result70[132]^and_result70[133]^and_result70[134]^and_result70[135]^and_result70[136]^and_result70[137]^and_result70[138]^and_result70[139]^and_result70[140]^and_result70[141]^and_result70[142]^and_result70[143]^and_result70[144]^and_result70[145]^and_result70[146]^and_result70[147]^and_result70[148]^and_result70[149]^and_result70[150]^and_result70[151]^and_result70[152]^and_result70[153]^and_result70[154]^and_result70[155]^and_result70[156]^and_result70[157]^and_result70[158]^and_result70[159]^and_result70[160]^and_result70[161]^and_result70[162]^and_result70[163]^and_result70[164]^and_result70[165]^and_result70[166]^and_result70[167]^and_result70[168]^and_result70[169]^and_result70[170]^and_result70[171]^and_result70[172]^and_result70[173]^and_result70[174]^and_result70[175]^and_result70[176]^and_result70[177]^and_result70[178]^and_result70[179]^and_result70[180]^and_result70[181]^and_result70[182]^and_result70[183]^and_result70[184]^and_result70[185]^and_result70[186]^and_result70[187]^and_result70[188]^and_result70[189]^and_result70[190]^and_result70[191]^and_result70[192]^and_result70[193]^and_result70[194]^and_result70[195]^and_result70[196]^and_result70[197]^and_result70[198]^and_result70[199]^and_result70[200]^and_result70[201]^and_result70[202]^and_result70[203]^and_result70[204]^and_result70[205]^and_result70[206]^and_result70[207]^and_result70[208]^and_result70[209]^and_result70[210]^and_result70[211]^and_result70[212]^and_result70[213]^and_result70[214]^and_result70[215]^and_result70[216]^and_result70[217]^and_result70[218]^and_result70[219]^and_result70[220]^and_result70[221]^and_result70[222]^and_result70[223]^and_result70[224]^and_result70[225]^and_result70[226]^and_result70[227]^and_result70[228]^and_result70[229]^and_result70[230]^and_result70[231]^and_result70[232]^and_result70[233]^and_result70[234]^and_result70[235]^and_result70[236]^and_result70[237]^and_result70[238]^and_result70[239]^and_result70[240]^and_result70[241]^and_result70[242]^and_result70[243]^and_result70[244]^and_result70[245]^and_result70[246]^and_result70[247]^and_result70[248]^and_result70[249]^and_result70[250]^and_result70[251]^and_result70[252]^and_result70[253]^and_result70[254];
assign key[71]=and_result71[0]^and_result71[1]^and_result71[2]^and_result71[3]^and_result71[4]^and_result71[5]^and_result71[6]^and_result71[7]^and_result71[8]^and_result71[9]^and_result71[10]^and_result71[11]^and_result71[12]^and_result71[13]^and_result71[14]^and_result71[15]^and_result71[16]^and_result71[17]^and_result71[18]^and_result71[19]^and_result71[20]^and_result71[21]^and_result71[22]^and_result71[23]^and_result71[24]^and_result71[25]^and_result71[26]^and_result71[27]^and_result71[28]^and_result71[29]^and_result71[30]^and_result71[31]^and_result71[32]^and_result71[33]^and_result71[34]^and_result71[35]^and_result71[36]^and_result71[37]^and_result71[38]^and_result71[39]^and_result71[40]^and_result71[41]^and_result71[42]^and_result71[43]^and_result71[44]^and_result71[45]^and_result71[46]^and_result71[47]^and_result71[48]^and_result71[49]^and_result71[50]^and_result71[51]^and_result71[52]^and_result71[53]^and_result71[54]^and_result71[55]^and_result71[56]^and_result71[57]^and_result71[58]^and_result71[59]^and_result71[60]^and_result71[61]^and_result71[62]^and_result71[63]^and_result71[64]^and_result71[65]^and_result71[66]^and_result71[67]^and_result71[68]^and_result71[69]^and_result71[70]^and_result71[71]^and_result71[72]^and_result71[73]^and_result71[74]^and_result71[75]^and_result71[76]^and_result71[77]^and_result71[78]^and_result71[79]^and_result71[80]^and_result71[81]^and_result71[82]^and_result71[83]^and_result71[84]^and_result71[85]^and_result71[86]^and_result71[87]^and_result71[88]^and_result71[89]^and_result71[90]^and_result71[91]^and_result71[92]^and_result71[93]^and_result71[94]^and_result71[95]^and_result71[96]^and_result71[97]^and_result71[98]^and_result71[99]^and_result71[100]^and_result71[101]^and_result71[102]^and_result71[103]^and_result71[104]^and_result71[105]^and_result71[106]^and_result71[107]^and_result71[108]^and_result71[109]^and_result71[110]^and_result71[111]^and_result71[112]^and_result71[113]^and_result71[114]^and_result71[115]^and_result71[116]^and_result71[117]^and_result71[118]^and_result71[119]^and_result71[120]^and_result71[121]^and_result71[122]^and_result71[123]^and_result71[124]^and_result71[125]^and_result71[126]^and_result71[127]^and_result71[128]^and_result71[129]^and_result71[130]^and_result71[131]^and_result71[132]^and_result71[133]^and_result71[134]^and_result71[135]^and_result71[136]^and_result71[137]^and_result71[138]^and_result71[139]^and_result71[140]^and_result71[141]^and_result71[142]^and_result71[143]^and_result71[144]^and_result71[145]^and_result71[146]^and_result71[147]^and_result71[148]^and_result71[149]^and_result71[150]^and_result71[151]^and_result71[152]^and_result71[153]^and_result71[154]^and_result71[155]^and_result71[156]^and_result71[157]^and_result71[158]^and_result71[159]^and_result71[160]^and_result71[161]^and_result71[162]^and_result71[163]^and_result71[164]^and_result71[165]^and_result71[166]^and_result71[167]^and_result71[168]^and_result71[169]^and_result71[170]^and_result71[171]^and_result71[172]^and_result71[173]^and_result71[174]^and_result71[175]^and_result71[176]^and_result71[177]^and_result71[178]^and_result71[179]^and_result71[180]^and_result71[181]^and_result71[182]^and_result71[183]^and_result71[184]^and_result71[185]^and_result71[186]^and_result71[187]^and_result71[188]^and_result71[189]^and_result71[190]^and_result71[191]^and_result71[192]^and_result71[193]^and_result71[194]^and_result71[195]^and_result71[196]^and_result71[197]^and_result71[198]^and_result71[199]^and_result71[200]^and_result71[201]^and_result71[202]^and_result71[203]^and_result71[204]^and_result71[205]^and_result71[206]^and_result71[207]^and_result71[208]^and_result71[209]^and_result71[210]^and_result71[211]^and_result71[212]^and_result71[213]^and_result71[214]^and_result71[215]^and_result71[216]^and_result71[217]^and_result71[218]^and_result71[219]^and_result71[220]^and_result71[221]^and_result71[222]^and_result71[223]^and_result71[224]^and_result71[225]^and_result71[226]^and_result71[227]^and_result71[228]^and_result71[229]^and_result71[230]^and_result71[231]^and_result71[232]^and_result71[233]^and_result71[234]^and_result71[235]^and_result71[236]^and_result71[237]^and_result71[238]^and_result71[239]^and_result71[240]^and_result71[241]^and_result71[242]^and_result71[243]^and_result71[244]^and_result71[245]^and_result71[246]^and_result71[247]^and_result71[248]^and_result71[249]^and_result71[250]^and_result71[251]^and_result71[252]^and_result71[253]^and_result71[254];
assign key[72]=and_result72[0]^and_result72[1]^and_result72[2]^and_result72[3]^and_result72[4]^and_result72[5]^and_result72[6]^and_result72[7]^and_result72[8]^and_result72[9]^and_result72[10]^and_result72[11]^and_result72[12]^and_result72[13]^and_result72[14]^and_result72[15]^and_result72[16]^and_result72[17]^and_result72[18]^and_result72[19]^and_result72[20]^and_result72[21]^and_result72[22]^and_result72[23]^and_result72[24]^and_result72[25]^and_result72[26]^and_result72[27]^and_result72[28]^and_result72[29]^and_result72[30]^and_result72[31]^and_result72[32]^and_result72[33]^and_result72[34]^and_result72[35]^and_result72[36]^and_result72[37]^and_result72[38]^and_result72[39]^and_result72[40]^and_result72[41]^and_result72[42]^and_result72[43]^and_result72[44]^and_result72[45]^and_result72[46]^and_result72[47]^and_result72[48]^and_result72[49]^and_result72[50]^and_result72[51]^and_result72[52]^and_result72[53]^and_result72[54]^and_result72[55]^and_result72[56]^and_result72[57]^and_result72[58]^and_result72[59]^and_result72[60]^and_result72[61]^and_result72[62]^and_result72[63]^and_result72[64]^and_result72[65]^and_result72[66]^and_result72[67]^and_result72[68]^and_result72[69]^and_result72[70]^and_result72[71]^and_result72[72]^and_result72[73]^and_result72[74]^and_result72[75]^and_result72[76]^and_result72[77]^and_result72[78]^and_result72[79]^and_result72[80]^and_result72[81]^and_result72[82]^and_result72[83]^and_result72[84]^and_result72[85]^and_result72[86]^and_result72[87]^and_result72[88]^and_result72[89]^and_result72[90]^and_result72[91]^and_result72[92]^and_result72[93]^and_result72[94]^and_result72[95]^and_result72[96]^and_result72[97]^and_result72[98]^and_result72[99]^and_result72[100]^and_result72[101]^and_result72[102]^and_result72[103]^and_result72[104]^and_result72[105]^and_result72[106]^and_result72[107]^and_result72[108]^and_result72[109]^and_result72[110]^and_result72[111]^and_result72[112]^and_result72[113]^and_result72[114]^and_result72[115]^and_result72[116]^and_result72[117]^and_result72[118]^and_result72[119]^and_result72[120]^and_result72[121]^and_result72[122]^and_result72[123]^and_result72[124]^and_result72[125]^and_result72[126]^and_result72[127]^and_result72[128]^and_result72[129]^and_result72[130]^and_result72[131]^and_result72[132]^and_result72[133]^and_result72[134]^and_result72[135]^and_result72[136]^and_result72[137]^and_result72[138]^and_result72[139]^and_result72[140]^and_result72[141]^and_result72[142]^and_result72[143]^and_result72[144]^and_result72[145]^and_result72[146]^and_result72[147]^and_result72[148]^and_result72[149]^and_result72[150]^and_result72[151]^and_result72[152]^and_result72[153]^and_result72[154]^and_result72[155]^and_result72[156]^and_result72[157]^and_result72[158]^and_result72[159]^and_result72[160]^and_result72[161]^and_result72[162]^and_result72[163]^and_result72[164]^and_result72[165]^and_result72[166]^and_result72[167]^and_result72[168]^and_result72[169]^and_result72[170]^and_result72[171]^and_result72[172]^and_result72[173]^and_result72[174]^and_result72[175]^and_result72[176]^and_result72[177]^and_result72[178]^and_result72[179]^and_result72[180]^and_result72[181]^and_result72[182]^and_result72[183]^and_result72[184]^and_result72[185]^and_result72[186]^and_result72[187]^and_result72[188]^and_result72[189]^and_result72[190]^and_result72[191]^and_result72[192]^and_result72[193]^and_result72[194]^and_result72[195]^and_result72[196]^and_result72[197]^and_result72[198]^and_result72[199]^and_result72[200]^and_result72[201]^and_result72[202]^and_result72[203]^and_result72[204]^and_result72[205]^and_result72[206]^and_result72[207]^and_result72[208]^and_result72[209]^and_result72[210]^and_result72[211]^and_result72[212]^and_result72[213]^and_result72[214]^and_result72[215]^and_result72[216]^and_result72[217]^and_result72[218]^and_result72[219]^and_result72[220]^and_result72[221]^and_result72[222]^and_result72[223]^and_result72[224]^and_result72[225]^and_result72[226]^and_result72[227]^and_result72[228]^and_result72[229]^and_result72[230]^and_result72[231]^and_result72[232]^and_result72[233]^and_result72[234]^and_result72[235]^and_result72[236]^and_result72[237]^and_result72[238]^and_result72[239]^and_result72[240]^and_result72[241]^and_result72[242]^and_result72[243]^and_result72[244]^and_result72[245]^and_result72[246]^and_result72[247]^and_result72[248]^and_result72[249]^and_result72[250]^and_result72[251]^and_result72[252]^and_result72[253]^and_result72[254];
assign key[73]=and_result73[0]^and_result73[1]^and_result73[2]^and_result73[3]^and_result73[4]^and_result73[5]^and_result73[6]^and_result73[7]^and_result73[8]^and_result73[9]^and_result73[10]^and_result73[11]^and_result73[12]^and_result73[13]^and_result73[14]^and_result73[15]^and_result73[16]^and_result73[17]^and_result73[18]^and_result73[19]^and_result73[20]^and_result73[21]^and_result73[22]^and_result73[23]^and_result73[24]^and_result73[25]^and_result73[26]^and_result73[27]^and_result73[28]^and_result73[29]^and_result73[30]^and_result73[31]^and_result73[32]^and_result73[33]^and_result73[34]^and_result73[35]^and_result73[36]^and_result73[37]^and_result73[38]^and_result73[39]^and_result73[40]^and_result73[41]^and_result73[42]^and_result73[43]^and_result73[44]^and_result73[45]^and_result73[46]^and_result73[47]^and_result73[48]^and_result73[49]^and_result73[50]^and_result73[51]^and_result73[52]^and_result73[53]^and_result73[54]^and_result73[55]^and_result73[56]^and_result73[57]^and_result73[58]^and_result73[59]^and_result73[60]^and_result73[61]^and_result73[62]^and_result73[63]^and_result73[64]^and_result73[65]^and_result73[66]^and_result73[67]^and_result73[68]^and_result73[69]^and_result73[70]^and_result73[71]^and_result73[72]^and_result73[73]^and_result73[74]^and_result73[75]^and_result73[76]^and_result73[77]^and_result73[78]^and_result73[79]^and_result73[80]^and_result73[81]^and_result73[82]^and_result73[83]^and_result73[84]^and_result73[85]^and_result73[86]^and_result73[87]^and_result73[88]^and_result73[89]^and_result73[90]^and_result73[91]^and_result73[92]^and_result73[93]^and_result73[94]^and_result73[95]^and_result73[96]^and_result73[97]^and_result73[98]^and_result73[99]^and_result73[100]^and_result73[101]^and_result73[102]^and_result73[103]^and_result73[104]^and_result73[105]^and_result73[106]^and_result73[107]^and_result73[108]^and_result73[109]^and_result73[110]^and_result73[111]^and_result73[112]^and_result73[113]^and_result73[114]^and_result73[115]^and_result73[116]^and_result73[117]^and_result73[118]^and_result73[119]^and_result73[120]^and_result73[121]^and_result73[122]^and_result73[123]^and_result73[124]^and_result73[125]^and_result73[126]^and_result73[127]^and_result73[128]^and_result73[129]^and_result73[130]^and_result73[131]^and_result73[132]^and_result73[133]^and_result73[134]^and_result73[135]^and_result73[136]^and_result73[137]^and_result73[138]^and_result73[139]^and_result73[140]^and_result73[141]^and_result73[142]^and_result73[143]^and_result73[144]^and_result73[145]^and_result73[146]^and_result73[147]^and_result73[148]^and_result73[149]^and_result73[150]^and_result73[151]^and_result73[152]^and_result73[153]^and_result73[154]^and_result73[155]^and_result73[156]^and_result73[157]^and_result73[158]^and_result73[159]^and_result73[160]^and_result73[161]^and_result73[162]^and_result73[163]^and_result73[164]^and_result73[165]^and_result73[166]^and_result73[167]^and_result73[168]^and_result73[169]^and_result73[170]^and_result73[171]^and_result73[172]^and_result73[173]^and_result73[174]^and_result73[175]^and_result73[176]^and_result73[177]^and_result73[178]^and_result73[179]^and_result73[180]^and_result73[181]^and_result73[182]^and_result73[183]^and_result73[184]^and_result73[185]^and_result73[186]^and_result73[187]^and_result73[188]^and_result73[189]^and_result73[190]^and_result73[191]^and_result73[192]^and_result73[193]^and_result73[194]^and_result73[195]^and_result73[196]^and_result73[197]^and_result73[198]^and_result73[199]^and_result73[200]^and_result73[201]^and_result73[202]^and_result73[203]^and_result73[204]^and_result73[205]^and_result73[206]^and_result73[207]^and_result73[208]^and_result73[209]^and_result73[210]^and_result73[211]^and_result73[212]^and_result73[213]^and_result73[214]^and_result73[215]^and_result73[216]^and_result73[217]^and_result73[218]^and_result73[219]^and_result73[220]^and_result73[221]^and_result73[222]^and_result73[223]^and_result73[224]^and_result73[225]^and_result73[226]^and_result73[227]^and_result73[228]^and_result73[229]^and_result73[230]^and_result73[231]^and_result73[232]^and_result73[233]^and_result73[234]^and_result73[235]^and_result73[236]^and_result73[237]^and_result73[238]^and_result73[239]^and_result73[240]^and_result73[241]^and_result73[242]^and_result73[243]^and_result73[244]^and_result73[245]^and_result73[246]^and_result73[247]^and_result73[248]^and_result73[249]^and_result73[250]^and_result73[251]^and_result73[252]^and_result73[253]^and_result73[254];
assign key[74]=and_result74[0]^and_result74[1]^and_result74[2]^and_result74[3]^and_result74[4]^and_result74[5]^and_result74[6]^and_result74[7]^and_result74[8]^and_result74[9]^and_result74[10]^and_result74[11]^and_result74[12]^and_result74[13]^and_result74[14]^and_result74[15]^and_result74[16]^and_result74[17]^and_result74[18]^and_result74[19]^and_result74[20]^and_result74[21]^and_result74[22]^and_result74[23]^and_result74[24]^and_result74[25]^and_result74[26]^and_result74[27]^and_result74[28]^and_result74[29]^and_result74[30]^and_result74[31]^and_result74[32]^and_result74[33]^and_result74[34]^and_result74[35]^and_result74[36]^and_result74[37]^and_result74[38]^and_result74[39]^and_result74[40]^and_result74[41]^and_result74[42]^and_result74[43]^and_result74[44]^and_result74[45]^and_result74[46]^and_result74[47]^and_result74[48]^and_result74[49]^and_result74[50]^and_result74[51]^and_result74[52]^and_result74[53]^and_result74[54]^and_result74[55]^and_result74[56]^and_result74[57]^and_result74[58]^and_result74[59]^and_result74[60]^and_result74[61]^and_result74[62]^and_result74[63]^and_result74[64]^and_result74[65]^and_result74[66]^and_result74[67]^and_result74[68]^and_result74[69]^and_result74[70]^and_result74[71]^and_result74[72]^and_result74[73]^and_result74[74]^and_result74[75]^and_result74[76]^and_result74[77]^and_result74[78]^and_result74[79]^and_result74[80]^and_result74[81]^and_result74[82]^and_result74[83]^and_result74[84]^and_result74[85]^and_result74[86]^and_result74[87]^and_result74[88]^and_result74[89]^and_result74[90]^and_result74[91]^and_result74[92]^and_result74[93]^and_result74[94]^and_result74[95]^and_result74[96]^and_result74[97]^and_result74[98]^and_result74[99]^and_result74[100]^and_result74[101]^and_result74[102]^and_result74[103]^and_result74[104]^and_result74[105]^and_result74[106]^and_result74[107]^and_result74[108]^and_result74[109]^and_result74[110]^and_result74[111]^and_result74[112]^and_result74[113]^and_result74[114]^and_result74[115]^and_result74[116]^and_result74[117]^and_result74[118]^and_result74[119]^and_result74[120]^and_result74[121]^and_result74[122]^and_result74[123]^and_result74[124]^and_result74[125]^and_result74[126]^and_result74[127]^and_result74[128]^and_result74[129]^and_result74[130]^and_result74[131]^and_result74[132]^and_result74[133]^and_result74[134]^and_result74[135]^and_result74[136]^and_result74[137]^and_result74[138]^and_result74[139]^and_result74[140]^and_result74[141]^and_result74[142]^and_result74[143]^and_result74[144]^and_result74[145]^and_result74[146]^and_result74[147]^and_result74[148]^and_result74[149]^and_result74[150]^and_result74[151]^and_result74[152]^and_result74[153]^and_result74[154]^and_result74[155]^and_result74[156]^and_result74[157]^and_result74[158]^and_result74[159]^and_result74[160]^and_result74[161]^and_result74[162]^and_result74[163]^and_result74[164]^and_result74[165]^and_result74[166]^and_result74[167]^and_result74[168]^and_result74[169]^and_result74[170]^and_result74[171]^and_result74[172]^and_result74[173]^and_result74[174]^and_result74[175]^and_result74[176]^and_result74[177]^and_result74[178]^and_result74[179]^and_result74[180]^and_result74[181]^and_result74[182]^and_result74[183]^and_result74[184]^and_result74[185]^and_result74[186]^and_result74[187]^and_result74[188]^and_result74[189]^and_result74[190]^and_result74[191]^and_result74[192]^and_result74[193]^and_result74[194]^and_result74[195]^and_result74[196]^and_result74[197]^and_result74[198]^and_result74[199]^and_result74[200]^and_result74[201]^and_result74[202]^and_result74[203]^and_result74[204]^and_result74[205]^and_result74[206]^and_result74[207]^and_result74[208]^and_result74[209]^and_result74[210]^and_result74[211]^and_result74[212]^and_result74[213]^and_result74[214]^and_result74[215]^and_result74[216]^and_result74[217]^and_result74[218]^and_result74[219]^and_result74[220]^and_result74[221]^and_result74[222]^and_result74[223]^and_result74[224]^and_result74[225]^and_result74[226]^and_result74[227]^and_result74[228]^and_result74[229]^and_result74[230]^and_result74[231]^and_result74[232]^and_result74[233]^and_result74[234]^and_result74[235]^and_result74[236]^and_result74[237]^and_result74[238]^and_result74[239]^and_result74[240]^and_result74[241]^and_result74[242]^and_result74[243]^and_result74[244]^and_result74[245]^and_result74[246]^and_result74[247]^and_result74[248]^and_result74[249]^and_result74[250]^and_result74[251]^and_result74[252]^and_result74[253]^and_result74[254];
assign key[75]=and_result75[0]^and_result75[1]^and_result75[2]^and_result75[3]^and_result75[4]^and_result75[5]^and_result75[6]^and_result75[7]^and_result75[8]^and_result75[9]^and_result75[10]^and_result75[11]^and_result75[12]^and_result75[13]^and_result75[14]^and_result75[15]^and_result75[16]^and_result75[17]^and_result75[18]^and_result75[19]^and_result75[20]^and_result75[21]^and_result75[22]^and_result75[23]^and_result75[24]^and_result75[25]^and_result75[26]^and_result75[27]^and_result75[28]^and_result75[29]^and_result75[30]^and_result75[31]^and_result75[32]^and_result75[33]^and_result75[34]^and_result75[35]^and_result75[36]^and_result75[37]^and_result75[38]^and_result75[39]^and_result75[40]^and_result75[41]^and_result75[42]^and_result75[43]^and_result75[44]^and_result75[45]^and_result75[46]^and_result75[47]^and_result75[48]^and_result75[49]^and_result75[50]^and_result75[51]^and_result75[52]^and_result75[53]^and_result75[54]^and_result75[55]^and_result75[56]^and_result75[57]^and_result75[58]^and_result75[59]^and_result75[60]^and_result75[61]^and_result75[62]^and_result75[63]^and_result75[64]^and_result75[65]^and_result75[66]^and_result75[67]^and_result75[68]^and_result75[69]^and_result75[70]^and_result75[71]^and_result75[72]^and_result75[73]^and_result75[74]^and_result75[75]^and_result75[76]^and_result75[77]^and_result75[78]^and_result75[79]^and_result75[80]^and_result75[81]^and_result75[82]^and_result75[83]^and_result75[84]^and_result75[85]^and_result75[86]^and_result75[87]^and_result75[88]^and_result75[89]^and_result75[90]^and_result75[91]^and_result75[92]^and_result75[93]^and_result75[94]^and_result75[95]^and_result75[96]^and_result75[97]^and_result75[98]^and_result75[99]^and_result75[100]^and_result75[101]^and_result75[102]^and_result75[103]^and_result75[104]^and_result75[105]^and_result75[106]^and_result75[107]^and_result75[108]^and_result75[109]^and_result75[110]^and_result75[111]^and_result75[112]^and_result75[113]^and_result75[114]^and_result75[115]^and_result75[116]^and_result75[117]^and_result75[118]^and_result75[119]^and_result75[120]^and_result75[121]^and_result75[122]^and_result75[123]^and_result75[124]^and_result75[125]^and_result75[126]^and_result75[127]^and_result75[128]^and_result75[129]^and_result75[130]^and_result75[131]^and_result75[132]^and_result75[133]^and_result75[134]^and_result75[135]^and_result75[136]^and_result75[137]^and_result75[138]^and_result75[139]^and_result75[140]^and_result75[141]^and_result75[142]^and_result75[143]^and_result75[144]^and_result75[145]^and_result75[146]^and_result75[147]^and_result75[148]^and_result75[149]^and_result75[150]^and_result75[151]^and_result75[152]^and_result75[153]^and_result75[154]^and_result75[155]^and_result75[156]^and_result75[157]^and_result75[158]^and_result75[159]^and_result75[160]^and_result75[161]^and_result75[162]^and_result75[163]^and_result75[164]^and_result75[165]^and_result75[166]^and_result75[167]^and_result75[168]^and_result75[169]^and_result75[170]^and_result75[171]^and_result75[172]^and_result75[173]^and_result75[174]^and_result75[175]^and_result75[176]^and_result75[177]^and_result75[178]^and_result75[179]^and_result75[180]^and_result75[181]^and_result75[182]^and_result75[183]^and_result75[184]^and_result75[185]^and_result75[186]^and_result75[187]^and_result75[188]^and_result75[189]^and_result75[190]^and_result75[191]^and_result75[192]^and_result75[193]^and_result75[194]^and_result75[195]^and_result75[196]^and_result75[197]^and_result75[198]^and_result75[199]^and_result75[200]^and_result75[201]^and_result75[202]^and_result75[203]^and_result75[204]^and_result75[205]^and_result75[206]^and_result75[207]^and_result75[208]^and_result75[209]^and_result75[210]^and_result75[211]^and_result75[212]^and_result75[213]^and_result75[214]^and_result75[215]^and_result75[216]^and_result75[217]^and_result75[218]^and_result75[219]^and_result75[220]^and_result75[221]^and_result75[222]^and_result75[223]^and_result75[224]^and_result75[225]^and_result75[226]^and_result75[227]^and_result75[228]^and_result75[229]^and_result75[230]^and_result75[231]^and_result75[232]^and_result75[233]^and_result75[234]^and_result75[235]^and_result75[236]^and_result75[237]^and_result75[238]^and_result75[239]^and_result75[240]^and_result75[241]^and_result75[242]^and_result75[243]^and_result75[244]^and_result75[245]^and_result75[246]^and_result75[247]^and_result75[248]^and_result75[249]^and_result75[250]^and_result75[251]^and_result75[252]^and_result75[253]^and_result75[254];
assign key[76]=and_result76[0]^and_result76[1]^and_result76[2]^and_result76[3]^and_result76[4]^and_result76[5]^and_result76[6]^and_result76[7]^and_result76[8]^and_result76[9]^and_result76[10]^and_result76[11]^and_result76[12]^and_result76[13]^and_result76[14]^and_result76[15]^and_result76[16]^and_result76[17]^and_result76[18]^and_result76[19]^and_result76[20]^and_result76[21]^and_result76[22]^and_result76[23]^and_result76[24]^and_result76[25]^and_result76[26]^and_result76[27]^and_result76[28]^and_result76[29]^and_result76[30]^and_result76[31]^and_result76[32]^and_result76[33]^and_result76[34]^and_result76[35]^and_result76[36]^and_result76[37]^and_result76[38]^and_result76[39]^and_result76[40]^and_result76[41]^and_result76[42]^and_result76[43]^and_result76[44]^and_result76[45]^and_result76[46]^and_result76[47]^and_result76[48]^and_result76[49]^and_result76[50]^and_result76[51]^and_result76[52]^and_result76[53]^and_result76[54]^and_result76[55]^and_result76[56]^and_result76[57]^and_result76[58]^and_result76[59]^and_result76[60]^and_result76[61]^and_result76[62]^and_result76[63]^and_result76[64]^and_result76[65]^and_result76[66]^and_result76[67]^and_result76[68]^and_result76[69]^and_result76[70]^and_result76[71]^and_result76[72]^and_result76[73]^and_result76[74]^and_result76[75]^and_result76[76]^and_result76[77]^and_result76[78]^and_result76[79]^and_result76[80]^and_result76[81]^and_result76[82]^and_result76[83]^and_result76[84]^and_result76[85]^and_result76[86]^and_result76[87]^and_result76[88]^and_result76[89]^and_result76[90]^and_result76[91]^and_result76[92]^and_result76[93]^and_result76[94]^and_result76[95]^and_result76[96]^and_result76[97]^and_result76[98]^and_result76[99]^and_result76[100]^and_result76[101]^and_result76[102]^and_result76[103]^and_result76[104]^and_result76[105]^and_result76[106]^and_result76[107]^and_result76[108]^and_result76[109]^and_result76[110]^and_result76[111]^and_result76[112]^and_result76[113]^and_result76[114]^and_result76[115]^and_result76[116]^and_result76[117]^and_result76[118]^and_result76[119]^and_result76[120]^and_result76[121]^and_result76[122]^and_result76[123]^and_result76[124]^and_result76[125]^and_result76[126]^and_result76[127]^and_result76[128]^and_result76[129]^and_result76[130]^and_result76[131]^and_result76[132]^and_result76[133]^and_result76[134]^and_result76[135]^and_result76[136]^and_result76[137]^and_result76[138]^and_result76[139]^and_result76[140]^and_result76[141]^and_result76[142]^and_result76[143]^and_result76[144]^and_result76[145]^and_result76[146]^and_result76[147]^and_result76[148]^and_result76[149]^and_result76[150]^and_result76[151]^and_result76[152]^and_result76[153]^and_result76[154]^and_result76[155]^and_result76[156]^and_result76[157]^and_result76[158]^and_result76[159]^and_result76[160]^and_result76[161]^and_result76[162]^and_result76[163]^and_result76[164]^and_result76[165]^and_result76[166]^and_result76[167]^and_result76[168]^and_result76[169]^and_result76[170]^and_result76[171]^and_result76[172]^and_result76[173]^and_result76[174]^and_result76[175]^and_result76[176]^and_result76[177]^and_result76[178]^and_result76[179]^and_result76[180]^and_result76[181]^and_result76[182]^and_result76[183]^and_result76[184]^and_result76[185]^and_result76[186]^and_result76[187]^and_result76[188]^and_result76[189]^and_result76[190]^and_result76[191]^and_result76[192]^and_result76[193]^and_result76[194]^and_result76[195]^and_result76[196]^and_result76[197]^and_result76[198]^and_result76[199]^and_result76[200]^and_result76[201]^and_result76[202]^and_result76[203]^and_result76[204]^and_result76[205]^and_result76[206]^and_result76[207]^and_result76[208]^and_result76[209]^and_result76[210]^and_result76[211]^and_result76[212]^and_result76[213]^and_result76[214]^and_result76[215]^and_result76[216]^and_result76[217]^and_result76[218]^and_result76[219]^and_result76[220]^and_result76[221]^and_result76[222]^and_result76[223]^and_result76[224]^and_result76[225]^and_result76[226]^and_result76[227]^and_result76[228]^and_result76[229]^and_result76[230]^and_result76[231]^and_result76[232]^and_result76[233]^and_result76[234]^and_result76[235]^and_result76[236]^and_result76[237]^and_result76[238]^and_result76[239]^and_result76[240]^and_result76[241]^and_result76[242]^and_result76[243]^and_result76[244]^and_result76[245]^and_result76[246]^and_result76[247]^and_result76[248]^and_result76[249]^and_result76[250]^and_result76[251]^and_result76[252]^and_result76[253]^and_result76[254];
assign key[77]=and_result77[0]^and_result77[1]^and_result77[2]^and_result77[3]^and_result77[4]^and_result77[5]^and_result77[6]^and_result77[7]^and_result77[8]^and_result77[9]^and_result77[10]^and_result77[11]^and_result77[12]^and_result77[13]^and_result77[14]^and_result77[15]^and_result77[16]^and_result77[17]^and_result77[18]^and_result77[19]^and_result77[20]^and_result77[21]^and_result77[22]^and_result77[23]^and_result77[24]^and_result77[25]^and_result77[26]^and_result77[27]^and_result77[28]^and_result77[29]^and_result77[30]^and_result77[31]^and_result77[32]^and_result77[33]^and_result77[34]^and_result77[35]^and_result77[36]^and_result77[37]^and_result77[38]^and_result77[39]^and_result77[40]^and_result77[41]^and_result77[42]^and_result77[43]^and_result77[44]^and_result77[45]^and_result77[46]^and_result77[47]^and_result77[48]^and_result77[49]^and_result77[50]^and_result77[51]^and_result77[52]^and_result77[53]^and_result77[54]^and_result77[55]^and_result77[56]^and_result77[57]^and_result77[58]^and_result77[59]^and_result77[60]^and_result77[61]^and_result77[62]^and_result77[63]^and_result77[64]^and_result77[65]^and_result77[66]^and_result77[67]^and_result77[68]^and_result77[69]^and_result77[70]^and_result77[71]^and_result77[72]^and_result77[73]^and_result77[74]^and_result77[75]^and_result77[76]^and_result77[77]^and_result77[78]^and_result77[79]^and_result77[80]^and_result77[81]^and_result77[82]^and_result77[83]^and_result77[84]^and_result77[85]^and_result77[86]^and_result77[87]^and_result77[88]^and_result77[89]^and_result77[90]^and_result77[91]^and_result77[92]^and_result77[93]^and_result77[94]^and_result77[95]^and_result77[96]^and_result77[97]^and_result77[98]^and_result77[99]^and_result77[100]^and_result77[101]^and_result77[102]^and_result77[103]^and_result77[104]^and_result77[105]^and_result77[106]^and_result77[107]^and_result77[108]^and_result77[109]^and_result77[110]^and_result77[111]^and_result77[112]^and_result77[113]^and_result77[114]^and_result77[115]^and_result77[116]^and_result77[117]^and_result77[118]^and_result77[119]^and_result77[120]^and_result77[121]^and_result77[122]^and_result77[123]^and_result77[124]^and_result77[125]^and_result77[126]^and_result77[127]^and_result77[128]^and_result77[129]^and_result77[130]^and_result77[131]^and_result77[132]^and_result77[133]^and_result77[134]^and_result77[135]^and_result77[136]^and_result77[137]^and_result77[138]^and_result77[139]^and_result77[140]^and_result77[141]^and_result77[142]^and_result77[143]^and_result77[144]^and_result77[145]^and_result77[146]^and_result77[147]^and_result77[148]^and_result77[149]^and_result77[150]^and_result77[151]^and_result77[152]^and_result77[153]^and_result77[154]^and_result77[155]^and_result77[156]^and_result77[157]^and_result77[158]^and_result77[159]^and_result77[160]^and_result77[161]^and_result77[162]^and_result77[163]^and_result77[164]^and_result77[165]^and_result77[166]^and_result77[167]^and_result77[168]^and_result77[169]^and_result77[170]^and_result77[171]^and_result77[172]^and_result77[173]^and_result77[174]^and_result77[175]^and_result77[176]^and_result77[177]^and_result77[178]^and_result77[179]^and_result77[180]^and_result77[181]^and_result77[182]^and_result77[183]^and_result77[184]^and_result77[185]^and_result77[186]^and_result77[187]^and_result77[188]^and_result77[189]^and_result77[190]^and_result77[191]^and_result77[192]^and_result77[193]^and_result77[194]^and_result77[195]^and_result77[196]^and_result77[197]^and_result77[198]^and_result77[199]^and_result77[200]^and_result77[201]^and_result77[202]^and_result77[203]^and_result77[204]^and_result77[205]^and_result77[206]^and_result77[207]^and_result77[208]^and_result77[209]^and_result77[210]^and_result77[211]^and_result77[212]^and_result77[213]^and_result77[214]^and_result77[215]^and_result77[216]^and_result77[217]^and_result77[218]^and_result77[219]^and_result77[220]^and_result77[221]^and_result77[222]^and_result77[223]^and_result77[224]^and_result77[225]^and_result77[226]^and_result77[227]^and_result77[228]^and_result77[229]^and_result77[230]^and_result77[231]^and_result77[232]^and_result77[233]^and_result77[234]^and_result77[235]^and_result77[236]^and_result77[237]^and_result77[238]^and_result77[239]^and_result77[240]^and_result77[241]^and_result77[242]^and_result77[243]^and_result77[244]^and_result77[245]^and_result77[246]^and_result77[247]^and_result77[248]^and_result77[249]^and_result77[250]^and_result77[251]^and_result77[252]^and_result77[253]^and_result77[254];
assign key[78]=and_result78[0]^and_result78[1]^and_result78[2]^and_result78[3]^and_result78[4]^and_result78[5]^and_result78[6]^and_result78[7]^and_result78[8]^and_result78[9]^and_result78[10]^and_result78[11]^and_result78[12]^and_result78[13]^and_result78[14]^and_result78[15]^and_result78[16]^and_result78[17]^and_result78[18]^and_result78[19]^and_result78[20]^and_result78[21]^and_result78[22]^and_result78[23]^and_result78[24]^and_result78[25]^and_result78[26]^and_result78[27]^and_result78[28]^and_result78[29]^and_result78[30]^and_result78[31]^and_result78[32]^and_result78[33]^and_result78[34]^and_result78[35]^and_result78[36]^and_result78[37]^and_result78[38]^and_result78[39]^and_result78[40]^and_result78[41]^and_result78[42]^and_result78[43]^and_result78[44]^and_result78[45]^and_result78[46]^and_result78[47]^and_result78[48]^and_result78[49]^and_result78[50]^and_result78[51]^and_result78[52]^and_result78[53]^and_result78[54]^and_result78[55]^and_result78[56]^and_result78[57]^and_result78[58]^and_result78[59]^and_result78[60]^and_result78[61]^and_result78[62]^and_result78[63]^and_result78[64]^and_result78[65]^and_result78[66]^and_result78[67]^and_result78[68]^and_result78[69]^and_result78[70]^and_result78[71]^and_result78[72]^and_result78[73]^and_result78[74]^and_result78[75]^and_result78[76]^and_result78[77]^and_result78[78]^and_result78[79]^and_result78[80]^and_result78[81]^and_result78[82]^and_result78[83]^and_result78[84]^and_result78[85]^and_result78[86]^and_result78[87]^and_result78[88]^and_result78[89]^and_result78[90]^and_result78[91]^and_result78[92]^and_result78[93]^and_result78[94]^and_result78[95]^and_result78[96]^and_result78[97]^and_result78[98]^and_result78[99]^and_result78[100]^and_result78[101]^and_result78[102]^and_result78[103]^and_result78[104]^and_result78[105]^and_result78[106]^and_result78[107]^and_result78[108]^and_result78[109]^and_result78[110]^and_result78[111]^and_result78[112]^and_result78[113]^and_result78[114]^and_result78[115]^and_result78[116]^and_result78[117]^and_result78[118]^and_result78[119]^and_result78[120]^and_result78[121]^and_result78[122]^and_result78[123]^and_result78[124]^and_result78[125]^and_result78[126]^and_result78[127]^and_result78[128]^and_result78[129]^and_result78[130]^and_result78[131]^and_result78[132]^and_result78[133]^and_result78[134]^and_result78[135]^and_result78[136]^and_result78[137]^and_result78[138]^and_result78[139]^and_result78[140]^and_result78[141]^and_result78[142]^and_result78[143]^and_result78[144]^and_result78[145]^and_result78[146]^and_result78[147]^and_result78[148]^and_result78[149]^and_result78[150]^and_result78[151]^and_result78[152]^and_result78[153]^and_result78[154]^and_result78[155]^and_result78[156]^and_result78[157]^and_result78[158]^and_result78[159]^and_result78[160]^and_result78[161]^and_result78[162]^and_result78[163]^and_result78[164]^and_result78[165]^and_result78[166]^and_result78[167]^and_result78[168]^and_result78[169]^and_result78[170]^and_result78[171]^and_result78[172]^and_result78[173]^and_result78[174]^and_result78[175]^and_result78[176]^and_result78[177]^and_result78[178]^and_result78[179]^and_result78[180]^and_result78[181]^and_result78[182]^and_result78[183]^and_result78[184]^and_result78[185]^and_result78[186]^and_result78[187]^and_result78[188]^and_result78[189]^and_result78[190]^and_result78[191]^and_result78[192]^and_result78[193]^and_result78[194]^and_result78[195]^and_result78[196]^and_result78[197]^and_result78[198]^and_result78[199]^and_result78[200]^and_result78[201]^and_result78[202]^and_result78[203]^and_result78[204]^and_result78[205]^and_result78[206]^and_result78[207]^and_result78[208]^and_result78[209]^and_result78[210]^and_result78[211]^and_result78[212]^and_result78[213]^and_result78[214]^and_result78[215]^and_result78[216]^and_result78[217]^and_result78[218]^and_result78[219]^and_result78[220]^and_result78[221]^and_result78[222]^and_result78[223]^and_result78[224]^and_result78[225]^and_result78[226]^and_result78[227]^and_result78[228]^and_result78[229]^and_result78[230]^and_result78[231]^and_result78[232]^and_result78[233]^and_result78[234]^and_result78[235]^and_result78[236]^and_result78[237]^and_result78[238]^and_result78[239]^and_result78[240]^and_result78[241]^and_result78[242]^and_result78[243]^and_result78[244]^and_result78[245]^and_result78[246]^and_result78[247]^and_result78[248]^and_result78[249]^and_result78[250]^and_result78[251]^and_result78[252]^and_result78[253]^and_result78[254];
assign key[79]=and_result79[0]^and_result79[1]^and_result79[2]^and_result79[3]^and_result79[4]^and_result79[5]^and_result79[6]^and_result79[7]^and_result79[8]^and_result79[9]^and_result79[10]^and_result79[11]^and_result79[12]^and_result79[13]^and_result79[14]^and_result79[15]^and_result79[16]^and_result79[17]^and_result79[18]^and_result79[19]^and_result79[20]^and_result79[21]^and_result79[22]^and_result79[23]^and_result79[24]^and_result79[25]^and_result79[26]^and_result79[27]^and_result79[28]^and_result79[29]^and_result79[30]^and_result79[31]^and_result79[32]^and_result79[33]^and_result79[34]^and_result79[35]^and_result79[36]^and_result79[37]^and_result79[38]^and_result79[39]^and_result79[40]^and_result79[41]^and_result79[42]^and_result79[43]^and_result79[44]^and_result79[45]^and_result79[46]^and_result79[47]^and_result79[48]^and_result79[49]^and_result79[50]^and_result79[51]^and_result79[52]^and_result79[53]^and_result79[54]^and_result79[55]^and_result79[56]^and_result79[57]^and_result79[58]^and_result79[59]^and_result79[60]^and_result79[61]^and_result79[62]^and_result79[63]^and_result79[64]^and_result79[65]^and_result79[66]^and_result79[67]^and_result79[68]^and_result79[69]^and_result79[70]^and_result79[71]^and_result79[72]^and_result79[73]^and_result79[74]^and_result79[75]^and_result79[76]^and_result79[77]^and_result79[78]^and_result79[79]^and_result79[80]^and_result79[81]^and_result79[82]^and_result79[83]^and_result79[84]^and_result79[85]^and_result79[86]^and_result79[87]^and_result79[88]^and_result79[89]^and_result79[90]^and_result79[91]^and_result79[92]^and_result79[93]^and_result79[94]^and_result79[95]^and_result79[96]^and_result79[97]^and_result79[98]^and_result79[99]^and_result79[100]^and_result79[101]^and_result79[102]^and_result79[103]^and_result79[104]^and_result79[105]^and_result79[106]^and_result79[107]^and_result79[108]^and_result79[109]^and_result79[110]^and_result79[111]^and_result79[112]^and_result79[113]^and_result79[114]^and_result79[115]^and_result79[116]^and_result79[117]^and_result79[118]^and_result79[119]^and_result79[120]^and_result79[121]^and_result79[122]^and_result79[123]^and_result79[124]^and_result79[125]^and_result79[126]^and_result79[127]^and_result79[128]^and_result79[129]^and_result79[130]^and_result79[131]^and_result79[132]^and_result79[133]^and_result79[134]^and_result79[135]^and_result79[136]^and_result79[137]^and_result79[138]^and_result79[139]^and_result79[140]^and_result79[141]^and_result79[142]^and_result79[143]^and_result79[144]^and_result79[145]^and_result79[146]^and_result79[147]^and_result79[148]^and_result79[149]^and_result79[150]^and_result79[151]^and_result79[152]^and_result79[153]^and_result79[154]^and_result79[155]^and_result79[156]^and_result79[157]^and_result79[158]^and_result79[159]^and_result79[160]^and_result79[161]^and_result79[162]^and_result79[163]^and_result79[164]^and_result79[165]^and_result79[166]^and_result79[167]^and_result79[168]^and_result79[169]^and_result79[170]^and_result79[171]^and_result79[172]^and_result79[173]^and_result79[174]^and_result79[175]^and_result79[176]^and_result79[177]^and_result79[178]^and_result79[179]^and_result79[180]^and_result79[181]^and_result79[182]^and_result79[183]^and_result79[184]^and_result79[185]^and_result79[186]^and_result79[187]^and_result79[188]^and_result79[189]^and_result79[190]^and_result79[191]^and_result79[192]^and_result79[193]^and_result79[194]^and_result79[195]^and_result79[196]^and_result79[197]^and_result79[198]^and_result79[199]^and_result79[200]^and_result79[201]^and_result79[202]^and_result79[203]^and_result79[204]^and_result79[205]^and_result79[206]^and_result79[207]^and_result79[208]^and_result79[209]^and_result79[210]^and_result79[211]^and_result79[212]^and_result79[213]^and_result79[214]^and_result79[215]^and_result79[216]^and_result79[217]^and_result79[218]^and_result79[219]^and_result79[220]^and_result79[221]^and_result79[222]^and_result79[223]^and_result79[224]^and_result79[225]^and_result79[226]^and_result79[227]^and_result79[228]^and_result79[229]^and_result79[230]^and_result79[231]^and_result79[232]^and_result79[233]^and_result79[234]^and_result79[235]^and_result79[236]^and_result79[237]^and_result79[238]^and_result79[239]^and_result79[240]^and_result79[241]^and_result79[242]^and_result79[243]^and_result79[244]^and_result79[245]^and_result79[246]^and_result79[247]^and_result79[248]^and_result79[249]^and_result79[250]^and_result79[251]^and_result79[252]^and_result79[253]^and_result79[254];
assign key[80]=and_result80[0]^and_result80[1]^and_result80[2]^and_result80[3]^and_result80[4]^and_result80[5]^and_result80[6]^and_result80[7]^and_result80[8]^and_result80[9]^and_result80[10]^and_result80[11]^and_result80[12]^and_result80[13]^and_result80[14]^and_result80[15]^and_result80[16]^and_result80[17]^and_result80[18]^and_result80[19]^and_result80[20]^and_result80[21]^and_result80[22]^and_result80[23]^and_result80[24]^and_result80[25]^and_result80[26]^and_result80[27]^and_result80[28]^and_result80[29]^and_result80[30]^and_result80[31]^and_result80[32]^and_result80[33]^and_result80[34]^and_result80[35]^and_result80[36]^and_result80[37]^and_result80[38]^and_result80[39]^and_result80[40]^and_result80[41]^and_result80[42]^and_result80[43]^and_result80[44]^and_result80[45]^and_result80[46]^and_result80[47]^and_result80[48]^and_result80[49]^and_result80[50]^and_result80[51]^and_result80[52]^and_result80[53]^and_result80[54]^and_result80[55]^and_result80[56]^and_result80[57]^and_result80[58]^and_result80[59]^and_result80[60]^and_result80[61]^and_result80[62]^and_result80[63]^and_result80[64]^and_result80[65]^and_result80[66]^and_result80[67]^and_result80[68]^and_result80[69]^and_result80[70]^and_result80[71]^and_result80[72]^and_result80[73]^and_result80[74]^and_result80[75]^and_result80[76]^and_result80[77]^and_result80[78]^and_result80[79]^and_result80[80]^and_result80[81]^and_result80[82]^and_result80[83]^and_result80[84]^and_result80[85]^and_result80[86]^and_result80[87]^and_result80[88]^and_result80[89]^and_result80[90]^and_result80[91]^and_result80[92]^and_result80[93]^and_result80[94]^and_result80[95]^and_result80[96]^and_result80[97]^and_result80[98]^and_result80[99]^and_result80[100]^and_result80[101]^and_result80[102]^and_result80[103]^and_result80[104]^and_result80[105]^and_result80[106]^and_result80[107]^and_result80[108]^and_result80[109]^and_result80[110]^and_result80[111]^and_result80[112]^and_result80[113]^and_result80[114]^and_result80[115]^and_result80[116]^and_result80[117]^and_result80[118]^and_result80[119]^and_result80[120]^and_result80[121]^and_result80[122]^and_result80[123]^and_result80[124]^and_result80[125]^and_result80[126]^and_result80[127]^and_result80[128]^and_result80[129]^and_result80[130]^and_result80[131]^and_result80[132]^and_result80[133]^and_result80[134]^and_result80[135]^and_result80[136]^and_result80[137]^and_result80[138]^and_result80[139]^and_result80[140]^and_result80[141]^and_result80[142]^and_result80[143]^and_result80[144]^and_result80[145]^and_result80[146]^and_result80[147]^and_result80[148]^and_result80[149]^and_result80[150]^and_result80[151]^and_result80[152]^and_result80[153]^and_result80[154]^and_result80[155]^and_result80[156]^and_result80[157]^and_result80[158]^and_result80[159]^and_result80[160]^and_result80[161]^and_result80[162]^and_result80[163]^and_result80[164]^and_result80[165]^and_result80[166]^and_result80[167]^and_result80[168]^and_result80[169]^and_result80[170]^and_result80[171]^and_result80[172]^and_result80[173]^and_result80[174]^and_result80[175]^and_result80[176]^and_result80[177]^and_result80[178]^and_result80[179]^and_result80[180]^and_result80[181]^and_result80[182]^and_result80[183]^and_result80[184]^and_result80[185]^and_result80[186]^and_result80[187]^and_result80[188]^and_result80[189]^and_result80[190]^and_result80[191]^and_result80[192]^and_result80[193]^and_result80[194]^and_result80[195]^and_result80[196]^and_result80[197]^and_result80[198]^and_result80[199]^and_result80[200]^and_result80[201]^and_result80[202]^and_result80[203]^and_result80[204]^and_result80[205]^and_result80[206]^and_result80[207]^and_result80[208]^and_result80[209]^and_result80[210]^and_result80[211]^and_result80[212]^and_result80[213]^and_result80[214]^and_result80[215]^and_result80[216]^and_result80[217]^and_result80[218]^and_result80[219]^and_result80[220]^and_result80[221]^and_result80[222]^and_result80[223]^and_result80[224]^and_result80[225]^and_result80[226]^and_result80[227]^and_result80[228]^and_result80[229]^and_result80[230]^and_result80[231]^and_result80[232]^and_result80[233]^and_result80[234]^and_result80[235]^and_result80[236]^and_result80[237]^and_result80[238]^and_result80[239]^and_result80[240]^and_result80[241]^and_result80[242]^and_result80[243]^and_result80[244]^and_result80[245]^and_result80[246]^and_result80[247]^and_result80[248]^and_result80[249]^and_result80[250]^and_result80[251]^and_result80[252]^and_result80[253]^and_result80[254];
assign key[81]=and_result81[0]^and_result81[1]^and_result81[2]^and_result81[3]^and_result81[4]^and_result81[5]^and_result81[6]^and_result81[7]^and_result81[8]^and_result81[9]^and_result81[10]^and_result81[11]^and_result81[12]^and_result81[13]^and_result81[14]^and_result81[15]^and_result81[16]^and_result81[17]^and_result81[18]^and_result81[19]^and_result81[20]^and_result81[21]^and_result81[22]^and_result81[23]^and_result81[24]^and_result81[25]^and_result81[26]^and_result81[27]^and_result81[28]^and_result81[29]^and_result81[30]^and_result81[31]^and_result81[32]^and_result81[33]^and_result81[34]^and_result81[35]^and_result81[36]^and_result81[37]^and_result81[38]^and_result81[39]^and_result81[40]^and_result81[41]^and_result81[42]^and_result81[43]^and_result81[44]^and_result81[45]^and_result81[46]^and_result81[47]^and_result81[48]^and_result81[49]^and_result81[50]^and_result81[51]^and_result81[52]^and_result81[53]^and_result81[54]^and_result81[55]^and_result81[56]^and_result81[57]^and_result81[58]^and_result81[59]^and_result81[60]^and_result81[61]^and_result81[62]^and_result81[63]^and_result81[64]^and_result81[65]^and_result81[66]^and_result81[67]^and_result81[68]^and_result81[69]^and_result81[70]^and_result81[71]^and_result81[72]^and_result81[73]^and_result81[74]^and_result81[75]^and_result81[76]^and_result81[77]^and_result81[78]^and_result81[79]^and_result81[80]^and_result81[81]^and_result81[82]^and_result81[83]^and_result81[84]^and_result81[85]^and_result81[86]^and_result81[87]^and_result81[88]^and_result81[89]^and_result81[90]^and_result81[91]^and_result81[92]^and_result81[93]^and_result81[94]^and_result81[95]^and_result81[96]^and_result81[97]^and_result81[98]^and_result81[99]^and_result81[100]^and_result81[101]^and_result81[102]^and_result81[103]^and_result81[104]^and_result81[105]^and_result81[106]^and_result81[107]^and_result81[108]^and_result81[109]^and_result81[110]^and_result81[111]^and_result81[112]^and_result81[113]^and_result81[114]^and_result81[115]^and_result81[116]^and_result81[117]^and_result81[118]^and_result81[119]^and_result81[120]^and_result81[121]^and_result81[122]^and_result81[123]^and_result81[124]^and_result81[125]^and_result81[126]^and_result81[127]^and_result81[128]^and_result81[129]^and_result81[130]^and_result81[131]^and_result81[132]^and_result81[133]^and_result81[134]^and_result81[135]^and_result81[136]^and_result81[137]^and_result81[138]^and_result81[139]^and_result81[140]^and_result81[141]^and_result81[142]^and_result81[143]^and_result81[144]^and_result81[145]^and_result81[146]^and_result81[147]^and_result81[148]^and_result81[149]^and_result81[150]^and_result81[151]^and_result81[152]^and_result81[153]^and_result81[154]^and_result81[155]^and_result81[156]^and_result81[157]^and_result81[158]^and_result81[159]^and_result81[160]^and_result81[161]^and_result81[162]^and_result81[163]^and_result81[164]^and_result81[165]^and_result81[166]^and_result81[167]^and_result81[168]^and_result81[169]^and_result81[170]^and_result81[171]^and_result81[172]^and_result81[173]^and_result81[174]^and_result81[175]^and_result81[176]^and_result81[177]^and_result81[178]^and_result81[179]^and_result81[180]^and_result81[181]^and_result81[182]^and_result81[183]^and_result81[184]^and_result81[185]^and_result81[186]^and_result81[187]^and_result81[188]^and_result81[189]^and_result81[190]^and_result81[191]^and_result81[192]^and_result81[193]^and_result81[194]^and_result81[195]^and_result81[196]^and_result81[197]^and_result81[198]^and_result81[199]^and_result81[200]^and_result81[201]^and_result81[202]^and_result81[203]^and_result81[204]^and_result81[205]^and_result81[206]^and_result81[207]^and_result81[208]^and_result81[209]^and_result81[210]^and_result81[211]^and_result81[212]^and_result81[213]^and_result81[214]^and_result81[215]^and_result81[216]^and_result81[217]^and_result81[218]^and_result81[219]^and_result81[220]^and_result81[221]^and_result81[222]^and_result81[223]^and_result81[224]^and_result81[225]^and_result81[226]^and_result81[227]^and_result81[228]^and_result81[229]^and_result81[230]^and_result81[231]^and_result81[232]^and_result81[233]^and_result81[234]^and_result81[235]^and_result81[236]^and_result81[237]^and_result81[238]^and_result81[239]^and_result81[240]^and_result81[241]^and_result81[242]^and_result81[243]^and_result81[244]^and_result81[245]^and_result81[246]^and_result81[247]^and_result81[248]^and_result81[249]^and_result81[250]^and_result81[251]^and_result81[252]^and_result81[253]^and_result81[254];
assign key[82]=and_result82[0]^and_result82[1]^and_result82[2]^and_result82[3]^and_result82[4]^and_result82[5]^and_result82[6]^and_result82[7]^and_result82[8]^and_result82[9]^and_result82[10]^and_result82[11]^and_result82[12]^and_result82[13]^and_result82[14]^and_result82[15]^and_result82[16]^and_result82[17]^and_result82[18]^and_result82[19]^and_result82[20]^and_result82[21]^and_result82[22]^and_result82[23]^and_result82[24]^and_result82[25]^and_result82[26]^and_result82[27]^and_result82[28]^and_result82[29]^and_result82[30]^and_result82[31]^and_result82[32]^and_result82[33]^and_result82[34]^and_result82[35]^and_result82[36]^and_result82[37]^and_result82[38]^and_result82[39]^and_result82[40]^and_result82[41]^and_result82[42]^and_result82[43]^and_result82[44]^and_result82[45]^and_result82[46]^and_result82[47]^and_result82[48]^and_result82[49]^and_result82[50]^and_result82[51]^and_result82[52]^and_result82[53]^and_result82[54]^and_result82[55]^and_result82[56]^and_result82[57]^and_result82[58]^and_result82[59]^and_result82[60]^and_result82[61]^and_result82[62]^and_result82[63]^and_result82[64]^and_result82[65]^and_result82[66]^and_result82[67]^and_result82[68]^and_result82[69]^and_result82[70]^and_result82[71]^and_result82[72]^and_result82[73]^and_result82[74]^and_result82[75]^and_result82[76]^and_result82[77]^and_result82[78]^and_result82[79]^and_result82[80]^and_result82[81]^and_result82[82]^and_result82[83]^and_result82[84]^and_result82[85]^and_result82[86]^and_result82[87]^and_result82[88]^and_result82[89]^and_result82[90]^and_result82[91]^and_result82[92]^and_result82[93]^and_result82[94]^and_result82[95]^and_result82[96]^and_result82[97]^and_result82[98]^and_result82[99]^and_result82[100]^and_result82[101]^and_result82[102]^and_result82[103]^and_result82[104]^and_result82[105]^and_result82[106]^and_result82[107]^and_result82[108]^and_result82[109]^and_result82[110]^and_result82[111]^and_result82[112]^and_result82[113]^and_result82[114]^and_result82[115]^and_result82[116]^and_result82[117]^and_result82[118]^and_result82[119]^and_result82[120]^and_result82[121]^and_result82[122]^and_result82[123]^and_result82[124]^and_result82[125]^and_result82[126]^and_result82[127]^and_result82[128]^and_result82[129]^and_result82[130]^and_result82[131]^and_result82[132]^and_result82[133]^and_result82[134]^and_result82[135]^and_result82[136]^and_result82[137]^and_result82[138]^and_result82[139]^and_result82[140]^and_result82[141]^and_result82[142]^and_result82[143]^and_result82[144]^and_result82[145]^and_result82[146]^and_result82[147]^and_result82[148]^and_result82[149]^and_result82[150]^and_result82[151]^and_result82[152]^and_result82[153]^and_result82[154]^and_result82[155]^and_result82[156]^and_result82[157]^and_result82[158]^and_result82[159]^and_result82[160]^and_result82[161]^and_result82[162]^and_result82[163]^and_result82[164]^and_result82[165]^and_result82[166]^and_result82[167]^and_result82[168]^and_result82[169]^and_result82[170]^and_result82[171]^and_result82[172]^and_result82[173]^and_result82[174]^and_result82[175]^and_result82[176]^and_result82[177]^and_result82[178]^and_result82[179]^and_result82[180]^and_result82[181]^and_result82[182]^and_result82[183]^and_result82[184]^and_result82[185]^and_result82[186]^and_result82[187]^and_result82[188]^and_result82[189]^and_result82[190]^and_result82[191]^and_result82[192]^and_result82[193]^and_result82[194]^and_result82[195]^and_result82[196]^and_result82[197]^and_result82[198]^and_result82[199]^and_result82[200]^and_result82[201]^and_result82[202]^and_result82[203]^and_result82[204]^and_result82[205]^and_result82[206]^and_result82[207]^and_result82[208]^and_result82[209]^and_result82[210]^and_result82[211]^and_result82[212]^and_result82[213]^and_result82[214]^and_result82[215]^and_result82[216]^and_result82[217]^and_result82[218]^and_result82[219]^and_result82[220]^and_result82[221]^and_result82[222]^and_result82[223]^and_result82[224]^and_result82[225]^and_result82[226]^and_result82[227]^and_result82[228]^and_result82[229]^and_result82[230]^and_result82[231]^and_result82[232]^and_result82[233]^and_result82[234]^and_result82[235]^and_result82[236]^and_result82[237]^and_result82[238]^and_result82[239]^and_result82[240]^and_result82[241]^and_result82[242]^and_result82[243]^and_result82[244]^and_result82[245]^and_result82[246]^and_result82[247]^and_result82[248]^and_result82[249]^and_result82[250]^and_result82[251]^and_result82[252]^and_result82[253]^and_result82[254];
assign key[83]=and_result83[0]^and_result83[1]^and_result83[2]^and_result83[3]^and_result83[4]^and_result83[5]^and_result83[6]^and_result83[7]^and_result83[8]^and_result83[9]^and_result83[10]^and_result83[11]^and_result83[12]^and_result83[13]^and_result83[14]^and_result83[15]^and_result83[16]^and_result83[17]^and_result83[18]^and_result83[19]^and_result83[20]^and_result83[21]^and_result83[22]^and_result83[23]^and_result83[24]^and_result83[25]^and_result83[26]^and_result83[27]^and_result83[28]^and_result83[29]^and_result83[30]^and_result83[31]^and_result83[32]^and_result83[33]^and_result83[34]^and_result83[35]^and_result83[36]^and_result83[37]^and_result83[38]^and_result83[39]^and_result83[40]^and_result83[41]^and_result83[42]^and_result83[43]^and_result83[44]^and_result83[45]^and_result83[46]^and_result83[47]^and_result83[48]^and_result83[49]^and_result83[50]^and_result83[51]^and_result83[52]^and_result83[53]^and_result83[54]^and_result83[55]^and_result83[56]^and_result83[57]^and_result83[58]^and_result83[59]^and_result83[60]^and_result83[61]^and_result83[62]^and_result83[63]^and_result83[64]^and_result83[65]^and_result83[66]^and_result83[67]^and_result83[68]^and_result83[69]^and_result83[70]^and_result83[71]^and_result83[72]^and_result83[73]^and_result83[74]^and_result83[75]^and_result83[76]^and_result83[77]^and_result83[78]^and_result83[79]^and_result83[80]^and_result83[81]^and_result83[82]^and_result83[83]^and_result83[84]^and_result83[85]^and_result83[86]^and_result83[87]^and_result83[88]^and_result83[89]^and_result83[90]^and_result83[91]^and_result83[92]^and_result83[93]^and_result83[94]^and_result83[95]^and_result83[96]^and_result83[97]^and_result83[98]^and_result83[99]^and_result83[100]^and_result83[101]^and_result83[102]^and_result83[103]^and_result83[104]^and_result83[105]^and_result83[106]^and_result83[107]^and_result83[108]^and_result83[109]^and_result83[110]^and_result83[111]^and_result83[112]^and_result83[113]^and_result83[114]^and_result83[115]^and_result83[116]^and_result83[117]^and_result83[118]^and_result83[119]^and_result83[120]^and_result83[121]^and_result83[122]^and_result83[123]^and_result83[124]^and_result83[125]^and_result83[126]^and_result83[127]^and_result83[128]^and_result83[129]^and_result83[130]^and_result83[131]^and_result83[132]^and_result83[133]^and_result83[134]^and_result83[135]^and_result83[136]^and_result83[137]^and_result83[138]^and_result83[139]^and_result83[140]^and_result83[141]^and_result83[142]^and_result83[143]^and_result83[144]^and_result83[145]^and_result83[146]^and_result83[147]^and_result83[148]^and_result83[149]^and_result83[150]^and_result83[151]^and_result83[152]^and_result83[153]^and_result83[154]^and_result83[155]^and_result83[156]^and_result83[157]^and_result83[158]^and_result83[159]^and_result83[160]^and_result83[161]^and_result83[162]^and_result83[163]^and_result83[164]^and_result83[165]^and_result83[166]^and_result83[167]^and_result83[168]^and_result83[169]^and_result83[170]^and_result83[171]^and_result83[172]^and_result83[173]^and_result83[174]^and_result83[175]^and_result83[176]^and_result83[177]^and_result83[178]^and_result83[179]^and_result83[180]^and_result83[181]^and_result83[182]^and_result83[183]^and_result83[184]^and_result83[185]^and_result83[186]^and_result83[187]^and_result83[188]^and_result83[189]^and_result83[190]^and_result83[191]^and_result83[192]^and_result83[193]^and_result83[194]^and_result83[195]^and_result83[196]^and_result83[197]^and_result83[198]^and_result83[199]^and_result83[200]^and_result83[201]^and_result83[202]^and_result83[203]^and_result83[204]^and_result83[205]^and_result83[206]^and_result83[207]^and_result83[208]^and_result83[209]^and_result83[210]^and_result83[211]^and_result83[212]^and_result83[213]^and_result83[214]^and_result83[215]^and_result83[216]^and_result83[217]^and_result83[218]^and_result83[219]^and_result83[220]^and_result83[221]^and_result83[222]^and_result83[223]^and_result83[224]^and_result83[225]^and_result83[226]^and_result83[227]^and_result83[228]^and_result83[229]^and_result83[230]^and_result83[231]^and_result83[232]^and_result83[233]^and_result83[234]^and_result83[235]^and_result83[236]^and_result83[237]^and_result83[238]^and_result83[239]^and_result83[240]^and_result83[241]^and_result83[242]^and_result83[243]^and_result83[244]^and_result83[245]^and_result83[246]^and_result83[247]^and_result83[248]^and_result83[249]^and_result83[250]^and_result83[251]^and_result83[252]^and_result83[253]^and_result83[254];
assign key[84]=and_result84[0]^and_result84[1]^and_result84[2]^and_result84[3]^and_result84[4]^and_result84[5]^and_result84[6]^and_result84[7]^and_result84[8]^and_result84[9]^and_result84[10]^and_result84[11]^and_result84[12]^and_result84[13]^and_result84[14]^and_result84[15]^and_result84[16]^and_result84[17]^and_result84[18]^and_result84[19]^and_result84[20]^and_result84[21]^and_result84[22]^and_result84[23]^and_result84[24]^and_result84[25]^and_result84[26]^and_result84[27]^and_result84[28]^and_result84[29]^and_result84[30]^and_result84[31]^and_result84[32]^and_result84[33]^and_result84[34]^and_result84[35]^and_result84[36]^and_result84[37]^and_result84[38]^and_result84[39]^and_result84[40]^and_result84[41]^and_result84[42]^and_result84[43]^and_result84[44]^and_result84[45]^and_result84[46]^and_result84[47]^and_result84[48]^and_result84[49]^and_result84[50]^and_result84[51]^and_result84[52]^and_result84[53]^and_result84[54]^and_result84[55]^and_result84[56]^and_result84[57]^and_result84[58]^and_result84[59]^and_result84[60]^and_result84[61]^and_result84[62]^and_result84[63]^and_result84[64]^and_result84[65]^and_result84[66]^and_result84[67]^and_result84[68]^and_result84[69]^and_result84[70]^and_result84[71]^and_result84[72]^and_result84[73]^and_result84[74]^and_result84[75]^and_result84[76]^and_result84[77]^and_result84[78]^and_result84[79]^and_result84[80]^and_result84[81]^and_result84[82]^and_result84[83]^and_result84[84]^and_result84[85]^and_result84[86]^and_result84[87]^and_result84[88]^and_result84[89]^and_result84[90]^and_result84[91]^and_result84[92]^and_result84[93]^and_result84[94]^and_result84[95]^and_result84[96]^and_result84[97]^and_result84[98]^and_result84[99]^and_result84[100]^and_result84[101]^and_result84[102]^and_result84[103]^and_result84[104]^and_result84[105]^and_result84[106]^and_result84[107]^and_result84[108]^and_result84[109]^and_result84[110]^and_result84[111]^and_result84[112]^and_result84[113]^and_result84[114]^and_result84[115]^and_result84[116]^and_result84[117]^and_result84[118]^and_result84[119]^and_result84[120]^and_result84[121]^and_result84[122]^and_result84[123]^and_result84[124]^and_result84[125]^and_result84[126]^and_result84[127]^and_result84[128]^and_result84[129]^and_result84[130]^and_result84[131]^and_result84[132]^and_result84[133]^and_result84[134]^and_result84[135]^and_result84[136]^and_result84[137]^and_result84[138]^and_result84[139]^and_result84[140]^and_result84[141]^and_result84[142]^and_result84[143]^and_result84[144]^and_result84[145]^and_result84[146]^and_result84[147]^and_result84[148]^and_result84[149]^and_result84[150]^and_result84[151]^and_result84[152]^and_result84[153]^and_result84[154]^and_result84[155]^and_result84[156]^and_result84[157]^and_result84[158]^and_result84[159]^and_result84[160]^and_result84[161]^and_result84[162]^and_result84[163]^and_result84[164]^and_result84[165]^and_result84[166]^and_result84[167]^and_result84[168]^and_result84[169]^and_result84[170]^and_result84[171]^and_result84[172]^and_result84[173]^and_result84[174]^and_result84[175]^and_result84[176]^and_result84[177]^and_result84[178]^and_result84[179]^and_result84[180]^and_result84[181]^and_result84[182]^and_result84[183]^and_result84[184]^and_result84[185]^and_result84[186]^and_result84[187]^and_result84[188]^and_result84[189]^and_result84[190]^and_result84[191]^and_result84[192]^and_result84[193]^and_result84[194]^and_result84[195]^and_result84[196]^and_result84[197]^and_result84[198]^and_result84[199]^and_result84[200]^and_result84[201]^and_result84[202]^and_result84[203]^and_result84[204]^and_result84[205]^and_result84[206]^and_result84[207]^and_result84[208]^and_result84[209]^and_result84[210]^and_result84[211]^and_result84[212]^and_result84[213]^and_result84[214]^and_result84[215]^and_result84[216]^and_result84[217]^and_result84[218]^and_result84[219]^and_result84[220]^and_result84[221]^and_result84[222]^and_result84[223]^and_result84[224]^and_result84[225]^and_result84[226]^and_result84[227]^and_result84[228]^and_result84[229]^and_result84[230]^and_result84[231]^and_result84[232]^and_result84[233]^and_result84[234]^and_result84[235]^and_result84[236]^and_result84[237]^and_result84[238]^and_result84[239]^and_result84[240]^and_result84[241]^and_result84[242]^and_result84[243]^and_result84[244]^and_result84[245]^and_result84[246]^and_result84[247]^and_result84[248]^and_result84[249]^and_result84[250]^and_result84[251]^and_result84[252]^and_result84[253]^and_result84[254];
assign key[85]=and_result85[0]^and_result85[1]^and_result85[2]^and_result85[3]^and_result85[4]^and_result85[5]^and_result85[6]^and_result85[7]^and_result85[8]^and_result85[9]^and_result85[10]^and_result85[11]^and_result85[12]^and_result85[13]^and_result85[14]^and_result85[15]^and_result85[16]^and_result85[17]^and_result85[18]^and_result85[19]^and_result85[20]^and_result85[21]^and_result85[22]^and_result85[23]^and_result85[24]^and_result85[25]^and_result85[26]^and_result85[27]^and_result85[28]^and_result85[29]^and_result85[30]^and_result85[31]^and_result85[32]^and_result85[33]^and_result85[34]^and_result85[35]^and_result85[36]^and_result85[37]^and_result85[38]^and_result85[39]^and_result85[40]^and_result85[41]^and_result85[42]^and_result85[43]^and_result85[44]^and_result85[45]^and_result85[46]^and_result85[47]^and_result85[48]^and_result85[49]^and_result85[50]^and_result85[51]^and_result85[52]^and_result85[53]^and_result85[54]^and_result85[55]^and_result85[56]^and_result85[57]^and_result85[58]^and_result85[59]^and_result85[60]^and_result85[61]^and_result85[62]^and_result85[63]^and_result85[64]^and_result85[65]^and_result85[66]^and_result85[67]^and_result85[68]^and_result85[69]^and_result85[70]^and_result85[71]^and_result85[72]^and_result85[73]^and_result85[74]^and_result85[75]^and_result85[76]^and_result85[77]^and_result85[78]^and_result85[79]^and_result85[80]^and_result85[81]^and_result85[82]^and_result85[83]^and_result85[84]^and_result85[85]^and_result85[86]^and_result85[87]^and_result85[88]^and_result85[89]^and_result85[90]^and_result85[91]^and_result85[92]^and_result85[93]^and_result85[94]^and_result85[95]^and_result85[96]^and_result85[97]^and_result85[98]^and_result85[99]^and_result85[100]^and_result85[101]^and_result85[102]^and_result85[103]^and_result85[104]^and_result85[105]^and_result85[106]^and_result85[107]^and_result85[108]^and_result85[109]^and_result85[110]^and_result85[111]^and_result85[112]^and_result85[113]^and_result85[114]^and_result85[115]^and_result85[116]^and_result85[117]^and_result85[118]^and_result85[119]^and_result85[120]^and_result85[121]^and_result85[122]^and_result85[123]^and_result85[124]^and_result85[125]^and_result85[126]^and_result85[127]^and_result85[128]^and_result85[129]^and_result85[130]^and_result85[131]^and_result85[132]^and_result85[133]^and_result85[134]^and_result85[135]^and_result85[136]^and_result85[137]^and_result85[138]^and_result85[139]^and_result85[140]^and_result85[141]^and_result85[142]^and_result85[143]^and_result85[144]^and_result85[145]^and_result85[146]^and_result85[147]^and_result85[148]^and_result85[149]^and_result85[150]^and_result85[151]^and_result85[152]^and_result85[153]^and_result85[154]^and_result85[155]^and_result85[156]^and_result85[157]^and_result85[158]^and_result85[159]^and_result85[160]^and_result85[161]^and_result85[162]^and_result85[163]^and_result85[164]^and_result85[165]^and_result85[166]^and_result85[167]^and_result85[168]^and_result85[169]^and_result85[170]^and_result85[171]^and_result85[172]^and_result85[173]^and_result85[174]^and_result85[175]^and_result85[176]^and_result85[177]^and_result85[178]^and_result85[179]^and_result85[180]^and_result85[181]^and_result85[182]^and_result85[183]^and_result85[184]^and_result85[185]^and_result85[186]^and_result85[187]^and_result85[188]^and_result85[189]^and_result85[190]^and_result85[191]^and_result85[192]^and_result85[193]^and_result85[194]^and_result85[195]^and_result85[196]^and_result85[197]^and_result85[198]^and_result85[199]^and_result85[200]^and_result85[201]^and_result85[202]^and_result85[203]^and_result85[204]^and_result85[205]^and_result85[206]^and_result85[207]^and_result85[208]^and_result85[209]^and_result85[210]^and_result85[211]^and_result85[212]^and_result85[213]^and_result85[214]^and_result85[215]^and_result85[216]^and_result85[217]^and_result85[218]^and_result85[219]^and_result85[220]^and_result85[221]^and_result85[222]^and_result85[223]^and_result85[224]^and_result85[225]^and_result85[226]^and_result85[227]^and_result85[228]^and_result85[229]^and_result85[230]^and_result85[231]^and_result85[232]^and_result85[233]^and_result85[234]^and_result85[235]^and_result85[236]^and_result85[237]^and_result85[238]^and_result85[239]^and_result85[240]^and_result85[241]^and_result85[242]^and_result85[243]^and_result85[244]^and_result85[245]^and_result85[246]^and_result85[247]^and_result85[248]^and_result85[249]^and_result85[250]^and_result85[251]^and_result85[252]^and_result85[253]^and_result85[254];
assign key[86]=and_result86[0]^and_result86[1]^and_result86[2]^and_result86[3]^and_result86[4]^and_result86[5]^and_result86[6]^and_result86[7]^and_result86[8]^and_result86[9]^and_result86[10]^and_result86[11]^and_result86[12]^and_result86[13]^and_result86[14]^and_result86[15]^and_result86[16]^and_result86[17]^and_result86[18]^and_result86[19]^and_result86[20]^and_result86[21]^and_result86[22]^and_result86[23]^and_result86[24]^and_result86[25]^and_result86[26]^and_result86[27]^and_result86[28]^and_result86[29]^and_result86[30]^and_result86[31]^and_result86[32]^and_result86[33]^and_result86[34]^and_result86[35]^and_result86[36]^and_result86[37]^and_result86[38]^and_result86[39]^and_result86[40]^and_result86[41]^and_result86[42]^and_result86[43]^and_result86[44]^and_result86[45]^and_result86[46]^and_result86[47]^and_result86[48]^and_result86[49]^and_result86[50]^and_result86[51]^and_result86[52]^and_result86[53]^and_result86[54]^and_result86[55]^and_result86[56]^and_result86[57]^and_result86[58]^and_result86[59]^and_result86[60]^and_result86[61]^and_result86[62]^and_result86[63]^and_result86[64]^and_result86[65]^and_result86[66]^and_result86[67]^and_result86[68]^and_result86[69]^and_result86[70]^and_result86[71]^and_result86[72]^and_result86[73]^and_result86[74]^and_result86[75]^and_result86[76]^and_result86[77]^and_result86[78]^and_result86[79]^and_result86[80]^and_result86[81]^and_result86[82]^and_result86[83]^and_result86[84]^and_result86[85]^and_result86[86]^and_result86[87]^and_result86[88]^and_result86[89]^and_result86[90]^and_result86[91]^and_result86[92]^and_result86[93]^and_result86[94]^and_result86[95]^and_result86[96]^and_result86[97]^and_result86[98]^and_result86[99]^and_result86[100]^and_result86[101]^and_result86[102]^and_result86[103]^and_result86[104]^and_result86[105]^and_result86[106]^and_result86[107]^and_result86[108]^and_result86[109]^and_result86[110]^and_result86[111]^and_result86[112]^and_result86[113]^and_result86[114]^and_result86[115]^and_result86[116]^and_result86[117]^and_result86[118]^and_result86[119]^and_result86[120]^and_result86[121]^and_result86[122]^and_result86[123]^and_result86[124]^and_result86[125]^and_result86[126]^and_result86[127]^and_result86[128]^and_result86[129]^and_result86[130]^and_result86[131]^and_result86[132]^and_result86[133]^and_result86[134]^and_result86[135]^and_result86[136]^and_result86[137]^and_result86[138]^and_result86[139]^and_result86[140]^and_result86[141]^and_result86[142]^and_result86[143]^and_result86[144]^and_result86[145]^and_result86[146]^and_result86[147]^and_result86[148]^and_result86[149]^and_result86[150]^and_result86[151]^and_result86[152]^and_result86[153]^and_result86[154]^and_result86[155]^and_result86[156]^and_result86[157]^and_result86[158]^and_result86[159]^and_result86[160]^and_result86[161]^and_result86[162]^and_result86[163]^and_result86[164]^and_result86[165]^and_result86[166]^and_result86[167]^and_result86[168]^and_result86[169]^and_result86[170]^and_result86[171]^and_result86[172]^and_result86[173]^and_result86[174]^and_result86[175]^and_result86[176]^and_result86[177]^and_result86[178]^and_result86[179]^and_result86[180]^and_result86[181]^and_result86[182]^and_result86[183]^and_result86[184]^and_result86[185]^and_result86[186]^and_result86[187]^and_result86[188]^and_result86[189]^and_result86[190]^and_result86[191]^and_result86[192]^and_result86[193]^and_result86[194]^and_result86[195]^and_result86[196]^and_result86[197]^and_result86[198]^and_result86[199]^and_result86[200]^and_result86[201]^and_result86[202]^and_result86[203]^and_result86[204]^and_result86[205]^and_result86[206]^and_result86[207]^and_result86[208]^and_result86[209]^and_result86[210]^and_result86[211]^and_result86[212]^and_result86[213]^and_result86[214]^and_result86[215]^and_result86[216]^and_result86[217]^and_result86[218]^and_result86[219]^and_result86[220]^and_result86[221]^and_result86[222]^and_result86[223]^and_result86[224]^and_result86[225]^and_result86[226]^and_result86[227]^and_result86[228]^and_result86[229]^and_result86[230]^and_result86[231]^and_result86[232]^and_result86[233]^and_result86[234]^and_result86[235]^and_result86[236]^and_result86[237]^and_result86[238]^and_result86[239]^and_result86[240]^and_result86[241]^and_result86[242]^and_result86[243]^and_result86[244]^and_result86[245]^and_result86[246]^and_result86[247]^and_result86[248]^and_result86[249]^and_result86[250]^and_result86[251]^and_result86[252]^and_result86[253]^and_result86[254];
assign key[87]=and_result87[0]^and_result87[1]^and_result87[2]^and_result87[3]^and_result87[4]^and_result87[5]^and_result87[6]^and_result87[7]^and_result87[8]^and_result87[9]^and_result87[10]^and_result87[11]^and_result87[12]^and_result87[13]^and_result87[14]^and_result87[15]^and_result87[16]^and_result87[17]^and_result87[18]^and_result87[19]^and_result87[20]^and_result87[21]^and_result87[22]^and_result87[23]^and_result87[24]^and_result87[25]^and_result87[26]^and_result87[27]^and_result87[28]^and_result87[29]^and_result87[30]^and_result87[31]^and_result87[32]^and_result87[33]^and_result87[34]^and_result87[35]^and_result87[36]^and_result87[37]^and_result87[38]^and_result87[39]^and_result87[40]^and_result87[41]^and_result87[42]^and_result87[43]^and_result87[44]^and_result87[45]^and_result87[46]^and_result87[47]^and_result87[48]^and_result87[49]^and_result87[50]^and_result87[51]^and_result87[52]^and_result87[53]^and_result87[54]^and_result87[55]^and_result87[56]^and_result87[57]^and_result87[58]^and_result87[59]^and_result87[60]^and_result87[61]^and_result87[62]^and_result87[63]^and_result87[64]^and_result87[65]^and_result87[66]^and_result87[67]^and_result87[68]^and_result87[69]^and_result87[70]^and_result87[71]^and_result87[72]^and_result87[73]^and_result87[74]^and_result87[75]^and_result87[76]^and_result87[77]^and_result87[78]^and_result87[79]^and_result87[80]^and_result87[81]^and_result87[82]^and_result87[83]^and_result87[84]^and_result87[85]^and_result87[86]^and_result87[87]^and_result87[88]^and_result87[89]^and_result87[90]^and_result87[91]^and_result87[92]^and_result87[93]^and_result87[94]^and_result87[95]^and_result87[96]^and_result87[97]^and_result87[98]^and_result87[99]^and_result87[100]^and_result87[101]^and_result87[102]^and_result87[103]^and_result87[104]^and_result87[105]^and_result87[106]^and_result87[107]^and_result87[108]^and_result87[109]^and_result87[110]^and_result87[111]^and_result87[112]^and_result87[113]^and_result87[114]^and_result87[115]^and_result87[116]^and_result87[117]^and_result87[118]^and_result87[119]^and_result87[120]^and_result87[121]^and_result87[122]^and_result87[123]^and_result87[124]^and_result87[125]^and_result87[126]^and_result87[127]^and_result87[128]^and_result87[129]^and_result87[130]^and_result87[131]^and_result87[132]^and_result87[133]^and_result87[134]^and_result87[135]^and_result87[136]^and_result87[137]^and_result87[138]^and_result87[139]^and_result87[140]^and_result87[141]^and_result87[142]^and_result87[143]^and_result87[144]^and_result87[145]^and_result87[146]^and_result87[147]^and_result87[148]^and_result87[149]^and_result87[150]^and_result87[151]^and_result87[152]^and_result87[153]^and_result87[154]^and_result87[155]^and_result87[156]^and_result87[157]^and_result87[158]^and_result87[159]^and_result87[160]^and_result87[161]^and_result87[162]^and_result87[163]^and_result87[164]^and_result87[165]^and_result87[166]^and_result87[167]^and_result87[168]^and_result87[169]^and_result87[170]^and_result87[171]^and_result87[172]^and_result87[173]^and_result87[174]^and_result87[175]^and_result87[176]^and_result87[177]^and_result87[178]^and_result87[179]^and_result87[180]^and_result87[181]^and_result87[182]^and_result87[183]^and_result87[184]^and_result87[185]^and_result87[186]^and_result87[187]^and_result87[188]^and_result87[189]^and_result87[190]^and_result87[191]^and_result87[192]^and_result87[193]^and_result87[194]^and_result87[195]^and_result87[196]^and_result87[197]^and_result87[198]^and_result87[199]^and_result87[200]^and_result87[201]^and_result87[202]^and_result87[203]^and_result87[204]^and_result87[205]^and_result87[206]^and_result87[207]^and_result87[208]^and_result87[209]^and_result87[210]^and_result87[211]^and_result87[212]^and_result87[213]^and_result87[214]^and_result87[215]^and_result87[216]^and_result87[217]^and_result87[218]^and_result87[219]^and_result87[220]^and_result87[221]^and_result87[222]^and_result87[223]^and_result87[224]^and_result87[225]^and_result87[226]^and_result87[227]^and_result87[228]^and_result87[229]^and_result87[230]^and_result87[231]^and_result87[232]^and_result87[233]^and_result87[234]^and_result87[235]^and_result87[236]^and_result87[237]^and_result87[238]^and_result87[239]^and_result87[240]^and_result87[241]^and_result87[242]^and_result87[243]^and_result87[244]^and_result87[245]^and_result87[246]^and_result87[247]^and_result87[248]^and_result87[249]^and_result87[250]^and_result87[251]^and_result87[252]^and_result87[253]^and_result87[254];
assign key[88]=and_result88[0]^and_result88[1]^and_result88[2]^and_result88[3]^and_result88[4]^and_result88[5]^and_result88[6]^and_result88[7]^and_result88[8]^and_result88[9]^and_result88[10]^and_result88[11]^and_result88[12]^and_result88[13]^and_result88[14]^and_result88[15]^and_result88[16]^and_result88[17]^and_result88[18]^and_result88[19]^and_result88[20]^and_result88[21]^and_result88[22]^and_result88[23]^and_result88[24]^and_result88[25]^and_result88[26]^and_result88[27]^and_result88[28]^and_result88[29]^and_result88[30]^and_result88[31]^and_result88[32]^and_result88[33]^and_result88[34]^and_result88[35]^and_result88[36]^and_result88[37]^and_result88[38]^and_result88[39]^and_result88[40]^and_result88[41]^and_result88[42]^and_result88[43]^and_result88[44]^and_result88[45]^and_result88[46]^and_result88[47]^and_result88[48]^and_result88[49]^and_result88[50]^and_result88[51]^and_result88[52]^and_result88[53]^and_result88[54]^and_result88[55]^and_result88[56]^and_result88[57]^and_result88[58]^and_result88[59]^and_result88[60]^and_result88[61]^and_result88[62]^and_result88[63]^and_result88[64]^and_result88[65]^and_result88[66]^and_result88[67]^and_result88[68]^and_result88[69]^and_result88[70]^and_result88[71]^and_result88[72]^and_result88[73]^and_result88[74]^and_result88[75]^and_result88[76]^and_result88[77]^and_result88[78]^and_result88[79]^and_result88[80]^and_result88[81]^and_result88[82]^and_result88[83]^and_result88[84]^and_result88[85]^and_result88[86]^and_result88[87]^and_result88[88]^and_result88[89]^and_result88[90]^and_result88[91]^and_result88[92]^and_result88[93]^and_result88[94]^and_result88[95]^and_result88[96]^and_result88[97]^and_result88[98]^and_result88[99]^and_result88[100]^and_result88[101]^and_result88[102]^and_result88[103]^and_result88[104]^and_result88[105]^and_result88[106]^and_result88[107]^and_result88[108]^and_result88[109]^and_result88[110]^and_result88[111]^and_result88[112]^and_result88[113]^and_result88[114]^and_result88[115]^and_result88[116]^and_result88[117]^and_result88[118]^and_result88[119]^and_result88[120]^and_result88[121]^and_result88[122]^and_result88[123]^and_result88[124]^and_result88[125]^and_result88[126]^and_result88[127]^and_result88[128]^and_result88[129]^and_result88[130]^and_result88[131]^and_result88[132]^and_result88[133]^and_result88[134]^and_result88[135]^and_result88[136]^and_result88[137]^and_result88[138]^and_result88[139]^and_result88[140]^and_result88[141]^and_result88[142]^and_result88[143]^and_result88[144]^and_result88[145]^and_result88[146]^and_result88[147]^and_result88[148]^and_result88[149]^and_result88[150]^and_result88[151]^and_result88[152]^and_result88[153]^and_result88[154]^and_result88[155]^and_result88[156]^and_result88[157]^and_result88[158]^and_result88[159]^and_result88[160]^and_result88[161]^and_result88[162]^and_result88[163]^and_result88[164]^and_result88[165]^and_result88[166]^and_result88[167]^and_result88[168]^and_result88[169]^and_result88[170]^and_result88[171]^and_result88[172]^and_result88[173]^and_result88[174]^and_result88[175]^and_result88[176]^and_result88[177]^and_result88[178]^and_result88[179]^and_result88[180]^and_result88[181]^and_result88[182]^and_result88[183]^and_result88[184]^and_result88[185]^and_result88[186]^and_result88[187]^and_result88[188]^and_result88[189]^and_result88[190]^and_result88[191]^and_result88[192]^and_result88[193]^and_result88[194]^and_result88[195]^and_result88[196]^and_result88[197]^and_result88[198]^and_result88[199]^and_result88[200]^and_result88[201]^and_result88[202]^and_result88[203]^and_result88[204]^and_result88[205]^and_result88[206]^and_result88[207]^and_result88[208]^and_result88[209]^and_result88[210]^and_result88[211]^and_result88[212]^and_result88[213]^and_result88[214]^and_result88[215]^and_result88[216]^and_result88[217]^and_result88[218]^and_result88[219]^and_result88[220]^and_result88[221]^and_result88[222]^and_result88[223]^and_result88[224]^and_result88[225]^and_result88[226]^and_result88[227]^and_result88[228]^and_result88[229]^and_result88[230]^and_result88[231]^and_result88[232]^and_result88[233]^and_result88[234]^and_result88[235]^and_result88[236]^and_result88[237]^and_result88[238]^and_result88[239]^and_result88[240]^and_result88[241]^and_result88[242]^and_result88[243]^and_result88[244]^and_result88[245]^and_result88[246]^and_result88[247]^and_result88[248]^and_result88[249]^and_result88[250]^and_result88[251]^and_result88[252]^and_result88[253]^and_result88[254];
assign key[89]=and_result89[0]^and_result89[1]^and_result89[2]^and_result89[3]^and_result89[4]^and_result89[5]^and_result89[6]^and_result89[7]^and_result89[8]^and_result89[9]^and_result89[10]^and_result89[11]^and_result89[12]^and_result89[13]^and_result89[14]^and_result89[15]^and_result89[16]^and_result89[17]^and_result89[18]^and_result89[19]^and_result89[20]^and_result89[21]^and_result89[22]^and_result89[23]^and_result89[24]^and_result89[25]^and_result89[26]^and_result89[27]^and_result89[28]^and_result89[29]^and_result89[30]^and_result89[31]^and_result89[32]^and_result89[33]^and_result89[34]^and_result89[35]^and_result89[36]^and_result89[37]^and_result89[38]^and_result89[39]^and_result89[40]^and_result89[41]^and_result89[42]^and_result89[43]^and_result89[44]^and_result89[45]^and_result89[46]^and_result89[47]^and_result89[48]^and_result89[49]^and_result89[50]^and_result89[51]^and_result89[52]^and_result89[53]^and_result89[54]^and_result89[55]^and_result89[56]^and_result89[57]^and_result89[58]^and_result89[59]^and_result89[60]^and_result89[61]^and_result89[62]^and_result89[63]^and_result89[64]^and_result89[65]^and_result89[66]^and_result89[67]^and_result89[68]^and_result89[69]^and_result89[70]^and_result89[71]^and_result89[72]^and_result89[73]^and_result89[74]^and_result89[75]^and_result89[76]^and_result89[77]^and_result89[78]^and_result89[79]^and_result89[80]^and_result89[81]^and_result89[82]^and_result89[83]^and_result89[84]^and_result89[85]^and_result89[86]^and_result89[87]^and_result89[88]^and_result89[89]^and_result89[90]^and_result89[91]^and_result89[92]^and_result89[93]^and_result89[94]^and_result89[95]^and_result89[96]^and_result89[97]^and_result89[98]^and_result89[99]^and_result89[100]^and_result89[101]^and_result89[102]^and_result89[103]^and_result89[104]^and_result89[105]^and_result89[106]^and_result89[107]^and_result89[108]^and_result89[109]^and_result89[110]^and_result89[111]^and_result89[112]^and_result89[113]^and_result89[114]^and_result89[115]^and_result89[116]^and_result89[117]^and_result89[118]^and_result89[119]^and_result89[120]^and_result89[121]^and_result89[122]^and_result89[123]^and_result89[124]^and_result89[125]^and_result89[126]^and_result89[127]^and_result89[128]^and_result89[129]^and_result89[130]^and_result89[131]^and_result89[132]^and_result89[133]^and_result89[134]^and_result89[135]^and_result89[136]^and_result89[137]^and_result89[138]^and_result89[139]^and_result89[140]^and_result89[141]^and_result89[142]^and_result89[143]^and_result89[144]^and_result89[145]^and_result89[146]^and_result89[147]^and_result89[148]^and_result89[149]^and_result89[150]^and_result89[151]^and_result89[152]^and_result89[153]^and_result89[154]^and_result89[155]^and_result89[156]^and_result89[157]^and_result89[158]^and_result89[159]^and_result89[160]^and_result89[161]^and_result89[162]^and_result89[163]^and_result89[164]^and_result89[165]^and_result89[166]^and_result89[167]^and_result89[168]^and_result89[169]^and_result89[170]^and_result89[171]^and_result89[172]^and_result89[173]^and_result89[174]^and_result89[175]^and_result89[176]^and_result89[177]^and_result89[178]^and_result89[179]^and_result89[180]^and_result89[181]^and_result89[182]^and_result89[183]^and_result89[184]^and_result89[185]^and_result89[186]^and_result89[187]^and_result89[188]^and_result89[189]^and_result89[190]^and_result89[191]^and_result89[192]^and_result89[193]^and_result89[194]^and_result89[195]^and_result89[196]^and_result89[197]^and_result89[198]^and_result89[199]^and_result89[200]^and_result89[201]^and_result89[202]^and_result89[203]^and_result89[204]^and_result89[205]^and_result89[206]^and_result89[207]^and_result89[208]^and_result89[209]^and_result89[210]^and_result89[211]^and_result89[212]^and_result89[213]^and_result89[214]^and_result89[215]^and_result89[216]^and_result89[217]^and_result89[218]^and_result89[219]^and_result89[220]^and_result89[221]^and_result89[222]^and_result89[223]^and_result89[224]^and_result89[225]^and_result89[226]^and_result89[227]^and_result89[228]^and_result89[229]^and_result89[230]^and_result89[231]^and_result89[232]^and_result89[233]^and_result89[234]^and_result89[235]^and_result89[236]^and_result89[237]^and_result89[238]^and_result89[239]^and_result89[240]^and_result89[241]^and_result89[242]^and_result89[243]^and_result89[244]^and_result89[245]^and_result89[246]^and_result89[247]^and_result89[248]^and_result89[249]^and_result89[250]^and_result89[251]^and_result89[252]^and_result89[253]^and_result89[254];
assign key[90]=and_result90[0]^and_result90[1]^and_result90[2]^and_result90[3]^and_result90[4]^and_result90[5]^and_result90[6]^and_result90[7]^and_result90[8]^and_result90[9]^and_result90[10]^and_result90[11]^and_result90[12]^and_result90[13]^and_result90[14]^and_result90[15]^and_result90[16]^and_result90[17]^and_result90[18]^and_result90[19]^and_result90[20]^and_result90[21]^and_result90[22]^and_result90[23]^and_result90[24]^and_result90[25]^and_result90[26]^and_result90[27]^and_result90[28]^and_result90[29]^and_result90[30]^and_result90[31]^and_result90[32]^and_result90[33]^and_result90[34]^and_result90[35]^and_result90[36]^and_result90[37]^and_result90[38]^and_result90[39]^and_result90[40]^and_result90[41]^and_result90[42]^and_result90[43]^and_result90[44]^and_result90[45]^and_result90[46]^and_result90[47]^and_result90[48]^and_result90[49]^and_result90[50]^and_result90[51]^and_result90[52]^and_result90[53]^and_result90[54]^and_result90[55]^and_result90[56]^and_result90[57]^and_result90[58]^and_result90[59]^and_result90[60]^and_result90[61]^and_result90[62]^and_result90[63]^and_result90[64]^and_result90[65]^and_result90[66]^and_result90[67]^and_result90[68]^and_result90[69]^and_result90[70]^and_result90[71]^and_result90[72]^and_result90[73]^and_result90[74]^and_result90[75]^and_result90[76]^and_result90[77]^and_result90[78]^and_result90[79]^and_result90[80]^and_result90[81]^and_result90[82]^and_result90[83]^and_result90[84]^and_result90[85]^and_result90[86]^and_result90[87]^and_result90[88]^and_result90[89]^and_result90[90]^and_result90[91]^and_result90[92]^and_result90[93]^and_result90[94]^and_result90[95]^and_result90[96]^and_result90[97]^and_result90[98]^and_result90[99]^and_result90[100]^and_result90[101]^and_result90[102]^and_result90[103]^and_result90[104]^and_result90[105]^and_result90[106]^and_result90[107]^and_result90[108]^and_result90[109]^and_result90[110]^and_result90[111]^and_result90[112]^and_result90[113]^and_result90[114]^and_result90[115]^and_result90[116]^and_result90[117]^and_result90[118]^and_result90[119]^and_result90[120]^and_result90[121]^and_result90[122]^and_result90[123]^and_result90[124]^and_result90[125]^and_result90[126]^and_result90[127]^and_result90[128]^and_result90[129]^and_result90[130]^and_result90[131]^and_result90[132]^and_result90[133]^and_result90[134]^and_result90[135]^and_result90[136]^and_result90[137]^and_result90[138]^and_result90[139]^and_result90[140]^and_result90[141]^and_result90[142]^and_result90[143]^and_result90[144]^and_result90[145]^and_result90[146]^and_result90[147]^and_result90[148]^and_result90[149]^and_result90[150]^and_result90[151]^and_result90[152]^and_result90[153]^and_result90[154]^and_result90[155]^and_result90[156]^and_result90[157]^and_result90[158]^and_result90[159]^and_result90[160]^and_result90[161]^and_result90[162]^and_result90[163]^and_result90[164]^and_result90[165]^and_result90[166]^and_result90[167]^and_result90[168]^and_result90[169]^and_result90[170]^and_result90[171]^and_result90[172]^and_result90[173]^and_result90[174]^and_result90[175]^and_result90[176]^and_result90[177]^and_result90[178]^and_result90[179]^and_result90[180]^and_result90[181]^and_result90[182]^and_result90[183]^and_result90[184]^and_result90[185]^and_result90[186]^and_result90[187]^and_result90[188]^and_result90[189]^and_result90[190]^and_result90[191]^and_result90[192]^and_result90[193]^and_result90[194]^and_result90[195]^and_result90[196]^and_result90[197]^and_result90[198]^and_result90[199]^and_result90[200]^and_result90[201]^and_result90[202]^and_result90[203]^and_result90[204]^and_result90[205]^and_result90[206]^and_result90[207]^and_result90[208]^and_result90[209]^and_result90[210]^and_result90[211]^and_result90[212]^and_result90[213]^and_result90[214]^and_result90[215]^and_result90[216]^and_result90[217]^and_result90[218]^and_result90[219]^and_result90[220]^and_result90[221]^and_result90[222]^and_result90[223]^and_result90[224]^and_result90[225]^and_result90[226]^and_result90[227]^and_result90[228]^and_result90[229]^and_result90[230]^and_result90[231]^and_result90[232]^and_result90[233]^and_result90[234]^and_result90[235]^and_result90[236]^and_result90[237]^and_result90[238]^and_result90[239]^and_result90[240]^and_result90[241]^and_result90[242]^and_result90[243]^and_result90[244]^and_result90[245]^and_result90[246]^and_result90[247]^and_result90[248]^and_result90[249]^and_result90[250]^and_result90[251]^and_result90[252]^and_result90[253]^and_result90[254];
assign key[91]=and_result91[0]^and_result91[1]^and_result91[2]^and_result91[3]^and_result91[4]^and_result91[5]^and_result91[6]^and_result91[7]^and_result91[8]^and_result91[9]^and_result91[10]^and_result91[11]^and_result91[12]^and_result91[13]^and_result91[14]^and_result91[15]^and_result91[16]^and_result91[17]^and_result91[18]^and_result91[19]^and_result91[20]^and_result91[21]^and_result91[22]^and_result91[23]^and_result91[24]^and_result91[25]^and_result91[26]^and_result91[27]^and_result91[28]^and_result91[29]^and_result91[30]^and_result91[31]^and_result91[32]^and_result91[33]^and_result91[34]^and_result91[35]^and_result91[36]^and_result91[37]^and_result91[38]^and_result91[39]^and_result91[40]^and_result91[41]^and_result91[42]^and_result91[43]^and_result91[44]^and_result91[45]^and_result91[46]^and_result91[47]^and_result91[48]^and_result91[49]^and_result91[50]^and_result91[51]^and_result91[52]^and_result91[53]^and_result91[54]^and_result91[55]^and_result91[56]^and_result91[57]^and_result91[58]^and_result91[59]^and_result91[60]^and_result91[61]^and_result91[62]^and_result91[63]^and_result91[64]^and_result91[65]^and_result91[66]^and_result91[67]^and_result91[68]^and_result91[69]^and_result91[70]^and_result91[71]^and_result91[72]^and_result91[73]^and_result91[74]^and_result91[75]^and_result91[76]^and_result91[77]^and_result91[78]^and_result91[79]^and_result91[80]^and_result91[81]^and_result91[82]^and_result91[83]^and_result91[84]^and_result91[85]^and_result91[86]^and_result91[87]^and_result91[88]^and_result91[89]^and_result91[90]^and_result91[91]^and_result91[92]^and_result91[93]^and_result91[94]^and_result91[95]^and_result91[96]^and_result91[97]^and_result91[98]^and_result91[99]^and_result91[100]^and_result91[101]^and_result91[102]^and_result91[103]^and_result91[104]^and_result91[105]^and_result91[106]^and_result91[107]^and_result91[108]^and_result91[109]^and_result91[110]^and_result91[111]^and_result91[112]^and_result91[113]^and_result91[114]^and_result91[115]^and_result91[116]^and_result91[117]^and_result91[118]^and_result91[119]^and_result91[120]^and_result91[121]^and_result91[122]^and_result91[123]^and_result91[124]^and_result91[125]^and_result91[126]^and_result91[127]^and_result91[128]^and_result91[129]^and_result91[130]^and_result91[131]^and_result91[132]^and_result91[133]^and_result91[134]^and_result91[135]^and_result91[136]^and_result91[137]^and_result91[138]^and_result91[139]^and_result91[140]^and_result91[141]^and_result91[142]^and_result91[143]^and_result91[144]^and_result91[145]^and_result91[146]^and_result91[147]^and_result91[148]^and_result91[149]^and_result91[150]^and_result91[151]^and_result91[152]^and_result91[153]^and_result91[154]^and_result91[155]^and_result91[156]^and_result91[157]^and_result91[158]^and_result91[159]^and_result91[160]^and_result91[161]^and_result91[162]^and_result91[163]^and_result91[164]^and_result91[165]^and_result91[166]^and_result91[167]^and_result91[168]^and_result91[169]^and_result91[170]^and_result91[171]^and_result91[172]^and_result91[173]^and_result91[174]^and_result91[175]^and_result91[176]^and_result91[177]^and_result91[178]^and_result91[179]^and_result91[180]^and_result91[181]^and_result91[182]^and_result91[183]^and_result91[184]^and_result91[185]^and_result91[186]^and_result91[187]^and_result91[188]^and_result91[189]^and_result91[190]^and_result91[191]^and_result91[192]^and_result91[193]^and_result91[194]^and_result91[195]^and_result91[196]^and_result91[197]^and_result91[198]^and_result91[199]^and_result91[200]^and_result91[201]^and_result91[202]^and_result91[203]^and_result91[204]^and_result91[205]^and_result91[206]^and_result91[207]^and_result91[208]^and_result91[209]^and_result91[210]^and_result91[211]^and_result91[212]^and_result91[213]^and_result91[214]^and_result91[215]^and_result91[216]^and_result91[217]^and_result91[218]^and_result91[219]^and_result91[220]^and_result91[221]^and_result91[222]^and_result91[223]^and_result91[224]^and_result91[225]^and_result91[226]^and_result91[227]^and_result91[228]^and_result91[229]^and_result91[230]^and_result91[231]^and_result91[232]^and_result91[233]^and_result91[234]^and_result91[235]^and_result91[236]^and_result91[237]^and_result91[238]^and_result91[239]^and_result91[240]^and_result91[241]^and_result91[242]^and_result91[243]^and_result91[244]^and_result91[245]^and_result91[246]^and_result91[247]^and_result91[248]^and_result91[249]^and_result91[250]^and_result91[251]^and_result91[252]^and_result91[253]^and_result91[254];
assign key[92]=and_result92[0]^and_result92[1]^and_result92[2]^and_result92[3]^and_result92[4]^and_result92[5]^and_result92[6]^and_result92[7]^and_result92[8]^and_result92[9]^and_result92[10]^and_result92[11]^and_result92[12]^and_result92[13]^and_result92[14]^and_result92[15]^and_result92[16]^and_result92[17]^and_result92[18]^and_result92[19]^and_result92[20]^and_result92[21]^and_result92[22]^and_result92[23]^and_result92[24]^and_result92[25]^and_result92[26]^and_result92[27]^and_result92[28]^and_result92[29]^and_result92[30]^and_result92[31]^and_result92[32]^and_result92[33]^and_result92[34]^and_result92[35]^and_result92[36]^and_result92[37]^and_result92[38]^and_result92[39]^and_result92[40]^and_result92[41]^and_result92[42]^and_result92[43]^and_result92[44]^and_result92[45]^and_result92[46]^and_result92[47]^and_result92[48]^and_result92[49]^and_result92[50]^and_result92[51]^and_result92[52]^and_result92[53]^and_result92[54]^and_result92[55]^and_result92[56]^and_result92[57]^and_result92[58]^and_result92[59]^and_result92[60]^and_result92[61]^and_result92[62]^and_result92[63]^and_result92[64]^and_result92[65]^and_result92[66]^and_result92[67]^and_result92[68]^and_result92[69]^and_result92[70]^and_result92[71]^and_result92[72]^and_result92[73]^and_result92[74]^and_result92[75]^and_result92[76]^and_result92[77]^and_result92[78]^and_result92[79]^and_result92[80]^and_result92[81]^and_result92[82]^and_result92[83]^and_result92[84]^and_result92[85]^and_result92[86]^and_result92[87]^and_result92[88]^and_result92[89]^and_result92[90]^and_result92[91]^and_result92[92]^and_result92[93]^and_result92[94]^and_result92[95]^and_result92[96]^and_result92[97]^and_result92[98]^and_result92[99]^and_result92[100]^and_result92[101]^and_result92[102]^and_result92[103]^and_result92[104]^and_result92[105]^and_result92[106]^and_result92[107]^and_result92[108]^and_result92[109]^and_result92[110]^and_result92[111]^and_result92[112]^and_result92[113]^and_result92[114]^and_result92[115]^and_result92[116]^and_result92[117]^and_result92[118]^and_result92[119]^and_result92[120]^and_result92[121]^and_result92[122]^and_result92[123]^and_result92[124]^and_result92[125]^and_result92[126]^and_result92[127]^and_result92[128]^and_result92[129]^and_result92[130]^and_result92[131]^and_result92[132]^and_result92[133]^and_result92[134]^and_result92[135]^and_result92[136]^and_result92[137]^and_result92[138]^and_result92[139]^and_result92[140]^and_result92[141]^and_result92[142]^and_result92[143]^and_result92[144]^and_result92[145]^and_result92[146]^and_result92[147]^and_result92[148]^and_result92[149]^and_result92[150]^and_result92[151]^and_result92[152]^and_result92[153]^and_result92[154]^and_result92[155]^and_result92[156]^and_result92[157]^and_result92[158]^and_result92[159]^and_result92[160]^and_result92[161]^and_result92[162]^and_result92[163]^and_result92[164]^and_result92[165]^and_result92[166]^and_result92[167]^and_result92[168]^and_result92[169]^and_result92[170]^and_result92[171]^and_result92[172]^and_result92[173]^and_result92[174]^and_result92[175]^and_result92[176]^and_result92[177]^and_result92[178]^and_result92[179]^and_result92[180]^and_result92[181]^and_result92[182]^and_result92[183]^and_result92[184]^and_result92[185]^and_result92[186]^and_result92[187]^and_result92[188]^and_result92[189]^and_result92[190]^and_result92[191]^and_result92[192]^and_result92[193]^and_result92[194]^and_result92[195]^and_result92[196]^and_result92[197]^and_result92[198]^and_result92[199]^and_result92[200]^and_result92[201]^and_result92[202]^and_result92[203]^and_result92[204]^and_result92[205]^and_result92[206]^and_result92[207]^and_result92[208]^and_result92[209]^and_result92[210]^and_result92[211]^and_result92[212]^and_result92[213]^and_result92[214]^and_result92[215]^and_result92[216]^and_result92[217]^and_result92[218]^and_result92[219]^and_result92[220]^and_result92[221]^and_result92[222]^and_result92[223]^and_result92[224]^and_result92[225]^and_result92[226]^and_result92[227]^and_result92[228]^and_result92[229]^and_result92[230]^and_result92[231]^and_result92[232]^and_result92[233]^and_result92[234]^and_result92[235]^and_result92[236]^and_result92[237]^and_result92[238]^and_result92[239]^and_result92[240]^and_result92[241]^and_result92[242]^and_result92[243]^and_result92[244]^and_result92[245]^and_result92[246]^and_result92[247]^and_result92[248]^and_result92[249]^and_result92[250]^and_result92[251]^and_result92[252]^and_result92[253]^and_result92[254];
assign key[93]=and_result93[0]^and_result93[1]^and_result93[2]^and_result93[3]^and_result93[4]^and_result93[5]^and_result93[6]^and_result93[7]^and_result93[8]^and_result93[9]^and_result93[10]^and_result93[11]^and_result93[12]^and_result93[13]^and_result93[14]^and_result93[15]^and_result93[16]^and_result93[17]^and_result93[18]^and_result93[19]^and_result93[20]^and_result93[21]^and_result93[22]^and_result93[23]^and_result93[24]^and_result93[25]^and_result93[26]^and_result93[27]^and_result93[28]^and_result93[29]^and_result93[30]^and_result93[31]^and_result93[32]^and_result93[33]^and_result93[34]^and_result93[35]^and_result93[36]^and_result93[37]^and_result93[38]^and_result93[39]^and_result93[40]^and_result93[41]^and_result93[42]^and_result93[43]^and_result93[44]^and_result93[45]^and_result93[46]^and_result93[47]^and_result93[48]^and_result93[49]^and_result93[50]^and_result93[51]^and_result93[52]^and_result93[53]^and_result93[54]^and_result93[55]^and_result93[56]^and_result93[57]^and_result93[58]^and_result93[59]^and_result93[60]^and_result93[61]^and_result93[62]^and_result93[63]^and_result93[64]^and_result93[65]^and_result93[66]^and_result93[67]^and_result93[68]^and_result93[69]^and_result93[70]^and_result93[71]^and_result93[72]^and_result93[73]^and_result93[74]^and_result93[75]^and_result93[76]^and_result93[77]^and_result93[78]^and_result93[79]^and_result93[80]^and_result93[81]^and_result93[82]^and_result93[83]^and_result93[84]^and_result93[85]^and_result93[86]^and_result93[87]^and_result93[88]^and_result93[89]^and_result93[90]^and_result93[91]^and_result93[92]^and_result93[93]^and_result93[94]^and_result93[95]^and_result93[96]^and_result93[97]^and_result93[98]^and_result93[99]^and_result93[100]^and_result93[101]^and_result93[102]^and_result93[103]^and_result93[104]^and_result93[105]^and_result93[106]^and_result93[107]^and_result93[108]^and_result93[109]^and_result93[110]^and_result93[111]^and_result93[112]^and_result93[113]^and_result93[114]^and_result93[115]^and_result93[116]^and_result93[117]^and_result93[118]^and_result93[119]^and_result93[120]^and_result93[121]^and_result93[122]^and_result93[123]^and_result93[124]^and_result93[125]^and_result93[126]^and_result93[127]^and_result93[128]^and_result93[129]^and_result93[130]^and_result93[131]^and_result93[132]^and_result93[133]^and_result93[134]^and_result93[135]^and_result93[136]^and_result93[137]^and_result93[138]^and_result93[139]^and_result93[140]^and_result93[141]^and_result93[142]^and_result93[143]^and_result93[144]^and_result93[145]^and_result93[146]^and_result93[147]^and_result93[148]^and_result93[149]^and_result93[150]^and_result93[151]^and_result93[152]^and_result93[153]^and_result93[154]^and_result93[155]^and_result93[156]^and_result93[157]^and_result93[158]^and_result93[159]^and_result93[160]^and_result93[161]^and_result93[162]^and_result93[163]^and_result93[164]^and_result93[165]^and_result93[166]^and_result93[167]^and_result93[168]^and_result93[169]^and_result93[170]^and_result93[171]^and_result93[172]^and_result93[173]^and_result93[174]^and_result93[175]^and_result93[176]^and_result93[177]^and_result93[178]^and_result93[179]^and_result93[180]^and_result93[181]^and_result93[182]^and_result93[183]^and_result93[184]^and_result93[185]^and_result93[186]^and_result93[187]^and_result93[188]^and_result93[189]^and_result93[190]^and_result93[191]^and_result93[192]^and_result93[193]^and_result93[194]^and_result93[195]^and_result93[196]^and_result93[197]^and_result93[198]^and_result93[199]^and_result93[200]^and_result93[201]^and_result93[202]^and_result93[203]^and_result93[204]^and_result93[205]^and_result93[206]^and_result93[207]^and_result93[208]^and_result93[209]^and_result93[210]^and_result93[211]^and_result93[212]^and_result93[213]^and_result93[214]^and_result93[215]^and_result93[216]^and_result93[217]^and_result93[218]^and_result93[219]^and_result93[220]^and_result93[221]^and_result93[222]^and_result93[223]^and_result93[224]^and_result93[225]^and_result93[226]^and_result93[227]^and_result93[228]^and_result93[229]^and_result93[230]^and_result93[231]^and_result93[232]^and_result93[233]^and_result93[234]^and_result93[235]^and_result93[236]^and_result93[237]^and_result93[238]^and_result93[239]^and_result93[240]^and_result93[241]^and_result93[242]^and_result93[243]^and_result93[244]^and_result93[245]^and_result93[246]^and_result93[247]^and_result93[248]^and_result93[249]^and_result93[250]^and_result93[251]^and_result93[252]^and_result93[253]^and_result93[254];
assign key[94]=and_result94[0]^and_result94[1]^and_result94[2]^and_result94[3]^and_result94[4]^and_result94[5]^and_result94[6]^and_result94[7]^and_result94[8]^and_result94[9]^and_result94[10]^and_result94[11]^and_result94[12]^and_result94[13]^and_result94[14]^and_result94[15]^and_result94[16]^and_result94[17]^and_result94[18]^and_result94[19]^and_result94[20]^and_result94[21]^and_result94[22]^and_result94[23]^and_result94[24]^and_result94[25]^and_result94[26]^and_result94[27]^and_result94[28]^and_result94[29]^and_result94[30]^and_result94[31]^and_result94[32]^and_result94[33]^and_result94[34]^and_result94[35]^and_result94[36]^and_result94[37]^and_result94[38]^and_result94[39]^and_result94[40]^and_result94[41]^and_result94[42]^and_result94[43]^and_result94[44]^and_result94[45]^and_result94[46]^and_result94[47]^and_result94[48]^and_result94[49]^and_result94[50]^and_result94[51]^and_result94[52]^and_result94[53]^and_result94[54]^and_result94[55]^and_result94[56]^and_result94[57]^and_result94[58]^and_result94[59]^and_result94[60]^and_result94[61]^and_result94[62]^and_result94[63]^and_result94[64]^and_result94[65]^and_result94[66]^and_result94[67]^and_result94[68]^and_result94[69]^and_result94[70]^and_result94[71]^and_result94[72]^and_result94[73]^and_result94[74]^and_result94[75]^and_result94[76]^and_result94[77]^and_result94[78]^and_result94[79]^and_result94[80]^and_result94[81]^and_result94[82]^and_result94[83]^and_result94[84]^and_result94[85]^and_result94[86]^and_result94[87]^and_result94[88]^and_result94[89]^and_result94[90]^and_result94[91]^and_result94[92]^and_result94[93]^and_result94[94]^and_result94[95]^and_result94[96]^and_result94[97]^and_result94[98]^and_result94[99]^and_result94[100]^and_result94[101]^and_result94[102]^and_result94[103]^and_result94[104]^and_result94[105]^and_result94[106]^and_result94[107]^and_result94[108]^and_result94[109]^and_result94[110]^and_result94[111]^and_result94[112]^and_result94[113]^and_result94[114]^and_result94[115]^and_result94[116]^and_result94[117]^and_result94[118]^and_result94[119]^and_result94[120]^and_result94[121]^and_result94[122]^and_result94[123]^and_result94[124]^and_result94[125]^and_result94[126]^and_result94[127]^and_result94[128]^and_result94[129]^and_result94[130]^and_result94[131]^and_result94[132]^and_result94[133]^and_result94[134]^and_result94[135]^and_result94[136]^and_result94[137]^and_result94[138]^and_result94[139]^and_result94[140]^and_result94[141]^and_result94[142]^and_result94[143]^and_result94[144]^and_result94[145]^and_result94[146]^and_result94[147]^and_result94[148]^and_result94[149]^and_result94[150]^and_result94[151]^and_result94[152]^and_result94[153]^and_result94[154]^and_result94[155]^and_result94[156]^and_result94[157]^and_result94[158]^and_result94[159]^and_result94[160]^and_result94[161]^and_result94[162]^and_result94[163]^and_result94[164]^and_result94[165]^and_result94[166]^and_result94[167]^and_result94[168]^and_result94[169]^and_result94[170]^and_result94[171]^and_result94[172]^and_result94[173]^and_result94[174]^and_result94[175]^and_result94[176]^and_result94[177]^and_result94[178]^and_result94[179]^and_result94[180]^and_result94[181]^and_result94[182]^and_result94[183]^and_result94[184]^and_result94[185]^and_result94[186]^and_result94[187]^and_result94[188]^and_result94[189]^and_result94[190]^and_result94[191]^and_result94[192]^and_result94[193]^and_result94[194]^and_result94[195]^and_result94[196]^and_result94[197]^and_result94[198]^and_result94[199]^and_result94[200]^and_result94[201]^and_result94[202]^and_result94[203]^and_result94[204]^and_result94[205]^and_result94[206]^and_result94[207]^and_result94[208]^and_result94[209]^and_result94[210]^and_result94[211]^and_result94[212]^and_result94[213]^and_result94[214]^and_result94[215]^and_result94[216]^and_result94[217]^and_result94[218]^and_result94[219]^and_result94[220]^and_result94[221]^and_result94[222]^and_result94[223]^and_result94[224]^and_result94[225]^and_result94[226]^and_result94[227]^and_result94[228]^and_result94[229]^and_result94[230]^and_result94[231]^and_result94[232]^and_result94[233]^and_result94[234]^and_result94[235]^and_result94[236]^and_result94[237]^and_result94[238]^and_result94[239]^and_result94[240]^and_result94[241]^and_result94[242]^and_result94[243]^and_result94[244]^and_result94[245]^and_result94[246]^and_result94[247]^and_result94[248]^and_result94[249]^and_result94[250]^and_result94[251]^and_result94[252]^and_result94[253]^and_result94[254];
assign key[95]=and_result95[0]^and_result95[1]^and_result95[2]^and_result95[3]^and_result95[4]^and_result95[5]^and_result95[6]^and_result95[7]^and_result95[8]^and_result95[9]^and_result95[10]^and_result95[11]^and_result95[12]^and_result95[13]^and_result95[14]^and_result95[15]^and_result95[16]^and_result95[17]^and_result95[18]^and_result95[19]^and_result95[20]^and_result95[21]^and_result95[22]^and_result95[23]^and_result95[24]^and_result95[25]^and_result95[26]^and_result95[27]^and_result95[28]^and_result95[29]^and_result95[30]^and_result95[31]^and_result95[32]^and_result95[33]^and_result95[34]^and_result95[35]^and_result95[36]^and_result95[37]^and_result95[38]^and_result95[39]^and_result95[40]^and_result95[41]^and_result95[42]^and_result95[43]^and_result95[44]^and_result95[45]^and_result95[46]^and_result95[47]^and_result95[48]^and_result95[49]^and_result95[50]^and_result95[51]^and_result95[52]^and_result95[53]^and_result95[54]^and_result95[55]^and_result95[56]^and_result95[57]^and_result95[58]^and_result95[59]^and_result95[60]^and_result95[61]^and_result95[62]^and_result95[63]^and_result95[64]^and_result95[65]^and_result95[66]^and_result95[67]^and_result95[68]^and_result95[69]^and_result95[70]^and_result95[71]^and_result95[72]^and_result95[73]^and_result95[74]^and_result95[75]^and_result95[76]^and_result95[77]^and_result95[78]^and_result95[79]^and_result95[80]^and_result95[81]^and_result95[82]^and_result95[83]^and_result95[84]^and_result95[85]^and_result95[86]^and_result95[87]^and_result95[88]^and_result95[89]^and_result95[90]^and_result95[91]^and_result95[92]^and_result95[93]^and_result95[94]^and_result95[95]^and_result95[96]^and_result95[97]^and_result95[98]^and_result95[99]^and_result95[100]^and_result95[101]^and_result95[102]^and_result95[103]^and_result95[104]^and_result95[105]^and_result95[106]^and_result95[107]^and_result95[108]^and_result95[109]^and_result95[110]^and_result95[111]^and_result95[112]^and_result95[113]^and_result95[114]^and_result95[115]^and_result95[116]^and_result95[117]^and_result95[118]^and_result95[119]^and_result95[120]^and_result95[121]^and_result95[122]^and_result95[123]^and_result95[124]^and_result95[125]^and_result95[126]^and_result95[127]^and_result95[128]^and_result95[129]^and_result95[130]^and_result95[131]^and_result95[132]^and_result95[133]^and_result95[134]^and_result95[135]^and_result95[136]^and_result95[137]^and_result95[138]^and_result95[139]^and_result95[140]^and_result95[141]^and_result95[142]^and_result95[143]^and_result95[144]^and_result95[145]^and_result95[146]^and_result95[147]^and_result95[148]^and_result95[149]^and_result95[150]^and_result95[151]^and_result95[152]^and_result95[153]^and_result95[154]^and_result95[155]^and_result95[156]^and_result95[157]^and_result95[158]^and_result95[159]^and_result95[160]^and_result95[161]^and_result95[162]^and_result95[163]^and_result95[164]^and_result95[165]^and_result95[166]^and_result95[167]^and_result95[168]^and_result95[169]^and_result95[170]^and_result95[171]^and_result95[172]^and_result95[173]^and_result95[174]^and_result95[175]^and_result95[176]^and_result95[177]^and_result95[178]^and_result95[179]^and_result95[180]^and_result95[181]^and_result95[182]^and_result95[183]^and_result95[184]^and_result95[185]^and_result95[186]^and_result95[187]^and_result95[188]^and_result95[189]^and_result95[190]^and_result95[191]^and_result95[192]^and_result95[193]^and_result95[194]^and_result95[195]^and_result95[196]^and_result95[197]^and_result95[198]^and_result95[199]^and_result95[200]^and_result95[201]^and_result95[202]^and_result95[203]^and_result95[204]^and_result95[205]^and_result95[206]^and_result95[207]^and_result95[208]^and_result95[209]^and_result95[210]^and_result95[211]^and_result95[212]^and_result95[213]^and_result95[214]^and_result95[215]^and_result95[216]^and_result95[217]^and_result95[218]^and_result95[219]^and_result95[220]^and_result95[221]^and_result95[222]^and_result95[223]^and_result95[224]^and_result95[225]^and_result95[226]^and_result95[227]^and_result95[228]^and_result95[229]^and_result95[230]^and_result95[231]^and_result95[232]^and_result95[233]^and_result95[234]^and_result95[235]^and_result95[236]^and_result95[237]^and_result95[238]^and_result95[239]^and_result95[240]^and_result95[241]^and_result95[242]^and_result95[243]^and_result95[244]^and_result95[245]^and_result95[246]^and_result95[247]^and_result95[248]^and_result95[249]^and_result95[250]^and_result95[251]^and_result95[252]^and_result95[253]^and_result95[254];
assign key[96]=and_result96[0]^and_result96[1]^and_result96[2]^and_result96[3]^and_result96[4]^and_result96[5]^and_result96[6]^and_result96[7]^and_result96[8]^and_result96[9]^and_result96[10]^and_result96[11]^and_result96[12]^and_result96[13]^and_result96[14]^and_result96[15]^and_result96[16]^and_result96[17]^and_result96[18]^and_result96[19]^and_result96[20]^and_result96[21]^and_result96[22]^and_result96[23]^and_result96[24]^and_result96[25]^and_result96[26]^and_result96[27]^and_result96[28]^and_result96[29]^and_result96[30]^and_result96[31]^and_result96[32]^and_result96[33]^and_result96[34]^and_result96[35]^and_result96[36]^and_result96[37]^and_result96[38]^and_result96[39]^and_result96[40]^and_result96[41]^and_result96[42]^and_result96[43]^and_result96[44]^and_result96[45]^and_result96[46]^and_result96[47]^and_result96[48]^and_result96[49]^and_result96[50]^and_result96[51]^and_result96[52]^and_result96[53]^and_result96[54]^and_result96[55]^and_result96[56]^and_result96[57]^and_result96[58]^and_result96[59]^and_result96[60]^and_result96[61]^and_result96[62]^and_result96[63]^and_result96[64]^and_result96[65]^and_result96[66]^and_result96[67]^and_result96[68]^and_result96[69]^and_result96[70]^and_result96[71]^and_result96[72]^and_result96[73]^and_result96[74]^and_result96[75]^and_result96[76]^and_result96[77]^and_result96[78]^and_result96[79]^and_result96[80]^and_result96[81]^and_result96[82]^and_result96[83]^and_result96[84]^and_result96[85]^and_result96[86]^and_result96[87]^and_result96[88]^and_result96[89]^and_result96[90]^and_result96[91]^and_result96[92]^and_result96[93]^and_result96[94]^and_result96[95]^and_result96[96]^and_result96[97]^and_result96[98]^and_result96[99]^and_result96[100]^and_result96[101]^and_result96[102]^and_result96[103]^and_result96[104]^and_result96[105]^and_result96[106]^and_result96[107]^and_result96[108]^and_result96[109]^and_result96[110]^and_result96[111]^and_result96[112]^and_result96[113]^and_result96[114]^and_result96[115]^and_result96[116]^and_result96[117]^and_result96[118]^and_result96[119]^and_result96[120]^and_result96[121]^and_result96[122]^and_result96[123]^and_result96[124]^and_result96[125]^and_result96[126]^and_result96[127]^and_result96[128]^and_result96[129]^and_result96[130]^and_result96[131]^and_result96[132]^and_result96[133]^and_result96[134]^and_result96[135]^and_result96[136]^and_result96[137]^and_result96[138]^and_result96[139]^and_result96[140]^and_result96[141]^and_result96[142]^and_result96[143]^and_result96[144]^and_result96[145]^and_result96[146]^and_result96[147]^and_result96[148]^and_result96[149]^and_result96[150]^and_result96[151]^and_result96[152]^and_result96[153]^and_result96[154]^and_result96[155]^and_result96[156]^and_result96[157]^and_result96[158]^and_result96[159]^and_result96[160]^and_result96[161]^and_result96[162]^and_result96[163]^and_result96[164]^and_result96[165]^and_result96[166]^and_result96[167]^and_result96[168]^and_result96[169]^and_result96[170]^and_result96[171]^and_result96[172]^and_result96[173]^and_result96[174]^and_result96[175]^and_result96[176]^and_result96[177]^and_result96[178]^and_result96[179]^and_result96[180]^and_result96[181]^and_result96[182]^and_result96[183]^and_result96[184]^and_result96[185]^and_result96[186]^and_result96[187]^and_result96[188]^and_result96[189]^and_result96[190]^and_result96[191]^and_result96[192]^and_result96[193]^and_result96[194]^and_result96[195]^and_result96[196]^and_result96[197]^and_result96[198]^and_result96[199]^and_result96[200]^and_result96[201]^and_result96[202]^and_result96[203]^and_result96[204]^and_result96[205]^and_result96[206]^and_result96[207]^and_result96[208]^and_result96[209]^and_result96[210]^and_result96[211]^and_result96[212]^and_result96[213]^and_result96[214]^and_result96[215]^and_result96[216]^and_result96[217]^and_result96[218]^and_result96[219]^and_result96[220]^and_result96[221]^and_result96[222]^and_result96[223]^and_result96[224]^and_result96[225]^and_result96[226]^and_result96[227]^and_result96[228]^and_result96[229]^and_result96[230]^and_result96[231]^and_result96[232]^and_result96[233]^and_result96[234]^and_result96[235]^and_result96[236]^and_result96[237]^and_result96[238]^and_result96[239]^and_result96[240]^and_result96[241]^and_result96[242]^and_result96[243]^and_result96[244]^and_result96[245]^and_result96[246]^and_result96[247]^and_result96[248]^and_result96[249]^and_result96[250]^and_result96[251]^and_result96[252]^and_result96[253]^and_result96[254];
assign key[97]=and_result97[0]^and_result97[1]^and_result97[2]^and_result97[3]^and_result97[4]^and_result97[5]^and_result97[6]^and_result97[7]^and_result97[8]^and_result97[9]^and_result97[10]^and_result97[11]^and_result97[12]^and_result97[13]^and_result97[14]^and_result97[15]^and_result97[16]^and_result97[17]^and_result97[18]^and_result97[19]^and_result97[20]^and_result97[21]^and_result97[22]^and_result97[23]^and_result97[24]^and_result97[25]^and_result97[26]^and_result97[27]^and_result97[28]^and_result97[29]^and_result97[30]^and_result97[31]^and_result97[32]^and_result97[33]^and_result97[34]^and_result97[35]^and_result97[36]^and_result97[37]^and_result97[38]^and_result97[39]^and_result97[40]^and_result97[41]^and_result97[42]^and_result97[43]^and_result97[44]^and_result97[45]^and_result97[46]^and_result97[47]^and_result97[48]^and_result97[49]^and_result97[50]^and_result97[51]^and_result97[52]^and_result97[53]^and_result97[54]^and_result97[55]^and_result97[56]^and_result97[57]^and_result97[58]^and_result97[59]^and_result97[60]^and_result97[61]^and_result97[62]^and_result97[63]^and_result97[64]^and_result97[65]^and_result97[66]^and_result97[67]^and_result97[68]^and_result97[69]^and_result97[70]^and_result97[71]^and_result97[72]^and_result97[73]^and_result97[74]^and_result97[75]^and_result97[76]^and_result97[77]^and_result97[78]^and_result97[79]^and_result97[80]^and_result97[81]^and_result97[82]^and_result97[83]^and_result97[84]^and_result97[85]^and_result97[86]^and_result97[87]^and_result97[88]^and_result97[89]^and_result97[90]^and_result97[91]^and_result97[92]^and_result97[93]^and_result97[94]^and_result97[95]^and_result97[96]^and_result97[97]^and_result97[98]^and_result97[99]^and_result97[100]^and_result97[101]^and_result97[102]^and_result97[103]^and_result97[104]^and_result97[105]^and_result97[106]^and_result97[107]^and_result97[108]^and_result97[109]^and_result97[110]^and_result97[111]^and_result97[112]^and_result97[113]^and_result97[114]^and_result97[115]^and_result97[116]^and_result97[117]^and_result97[118]^and_result97[119]^and_result97[120]^and_result97[121]^and_result97[122]^and_result97[123]^and_result97[124]^and_result97[125]^and_result97[126]^and_result97[127]^and_result97[128]^and_result97[129]^and_result97[130]^and_result97[131]^and_result97[132]^and_result97[133]^and_result97[134]^and_result97[135]^and_result97[136]^and_result97[137]^and_result97[138]^and_result97[139]^and_result97[140]^and_result97[141]^and_result97[142]^and_result97[143]^and_result97[144]^and_result97[145]^and_result97[146]^and_result97[147]^and_result97[148]^and_result97[149]^and_result97[150]^and_result97[151]^and_result97[152]^and_result97[153]^and_result97[154]^and_result97[155]^and_result97[156]^and_result97[157]^and_result97[158]^and_result97[159]^and_result97[160]^and_result97[161]^and_result97[162]^and_result97[163]^and_result97[164]^and_result97[165]^and_result97[166]^and_result97[167]^and_result97[168]^and_result97[169]^and_result97[170]^and_result97[171]^and_result97[172]^and_result97[173]^and_result97[174]^and_result97[175]^and_result97[176]^and_result97[177]^and_result97[178]^and_result97[179]^and_result97[180]^and_result97[181]^and_result97[182]^and_result97[183]^and_result97[184]^and_result97[185]^and_result97[186]^and_result97[187]^and_result97[188]^and_result97[189]^and_result97[190]^and_result97[191]^and_result97[192]^and_result97[193]^and_result97[194]^and_result97[195]^and_result97[196]^and_result97[197]^and_result97[198]^and_result97[199]^and_result97[200]^and_result97[201]^and_result97[202]^and_result97[203]^and_result97[204]^and_result97[205]^and_result97[206]^and_result97[207]^and_result97[208]^and_result97[209]^and_result97[210]^and_result97[211]^and_result97[212]^and_result97[213]^and_result97[214]^and_result97[215]^and_result97[216]^and_result97[217]^and_result97[218]^and_result97[219]^and_result97[220]^and_result97[221]^and_result97[222]^and_result97[223]^and_result97[224]^and_result97[225]^and_result97[226]^and_result97[227]^and_result97[228]^and_result97[229]^and_result97[230]^and_result97[231]^and_result97[232]^and_result97[233]^and_result97[234]^and_result97[235]^and_result97[236]^and_result97[237]^and_result97[238]^and_result97[239]^and_result97[240]^and_result97[241]^and_result97[242]^and_result97[243]^and_result97[244]^and_result97[245]^and_result97[246]^and_result97[247]^and_result97[248]^and_result97[249]^and_result97[250]^and_result97[251]^and_result97[252]^and_result97[253]^and_result97[254];
assign key[98]=and_result98[0]^and_result98[1]^and_result98[2]^and_result98[3]^and_result98[4]^and_result98[5]^and_result98[6]^and_result98[7]^and_result98[8]^and_result98[9]^and_result98[10]^and_result98[11]^and_result98[12]^and_result98[13]^and_result98[14]^and_result98[15]^and_result98[16]^and_result98[17]^and_result98[18]^and_result98[19]^and_result98[20]^and_result98[21]^and_result98[22]^and_result98[23]^and_result98[24]^and_result98[25]^and_result98[26]^and_result98[27]^and_result98[28]^and_result98[29]^and_result98[30]^and_result98[31]^and_result98[32]^and_result98[33]^and_result98[34]^and_result98[35]^and_result98[36]^and_result98[37]^and_result98[38]^and_result98[39]^and_result98[40]^and_result98[41]^and_result98[42]^and_result98[43]^and_result98[44]^and_result98[45]^and_result98[46]^and_result98[47]^and_result98[48]^and_result98[49]^and_result98[50]^and_result98[51]^and_result98[52]^and_result98[53]^and_result98[54]^and_result98[55]^and_result98[56]^and_result98[57]^and_result98[58]^and_result98[59]^and_result98[60]^and_result98[61]^and_result98[62]^and_result98[63]^and_result98[64]^and_result98[65]^and_result98[66]^and_result98[67]^and_result98[68]^and_result98[69]^and_result98[70]^and_result98[71]^and_result98[72]^and_result98[73]^and_result98[74]^and_result98[75]^and_result98[76]^and_result98[77]^and_result98[78]^and_result98[79]^and_result98[80]^and_result98[81]^and_result98[82]^and_result98[83]^and_result98[84]^and_result98[85]^and_result98[86]^and_result98[87]^and_result98[88]^and_result98[89]^and_result98[90]^and_result98[91]^and_result98[92]^and_result98[93]^and_result98[94]^and_result98[95]^and_result98[96]^and_result98[97]^and_result98[98]^and_result98[99]^and_result98[100]^and_result98[101]^and_result98[102]^and_result98[103]^and_result98[104]^and_result98[105]^and_result98[106]^and_result98[107]^and_result98[108]^and_result98[109]^and_result98[110]^and_result98[111]^and_result98[112]^and_result98[113]^and_result98[114]^and_result98[115]^and_result98[116]^and_result98[117]^and_result98[118]^and_result98[119]^and_result98[120]^and_result98[121]^and_result98[122]^and_result98[123]^and_result98[124]^and_result98[125]^and_result98[126]^and_result98[127]^and_result98[128]^and_result98[129]^and_result98[130]^and_result98[131]^and_result98[132]^and_result98[133]^and_result98[134]^and_result98[135]^and_result98[136]^and_result98[137]^and_result98[138]^and_result98[139]^and_result98[140]^and_result98[141]^and_result98[142]^and_result98[143]^and_result98[144]^and_result98[145]^and_result98[146]^and_result98[147]^and_result98[148]^and_result98[149]^and_result98[150]^and_result98[151]^and_result98[152]^and_result98[153]^and_result98[154]^and_result98[155]^and_result98[156]^and_result98[157]^and_result98[158]^and_result98[159]^and_result98[160]^and_result98[161]^and_result98[162]^and_result98[163]^and_result98[164]^and_result98[165]^and_result98[166]^and_result98[167]^and_result98[168]^and_result98[169]^and_result98[170]^and_result98[171]^and_result98[172]^and_result98[173]^and_result98[174]^and_result98[175]^and_result98[176]^and_result98[177]^and_result98[178]^and_result98[179]^and_result98[180]^and_result98[181]^and_result98[182]^and_result98[183]^and_result98[184]^and_result98[185]^and_result98[186]^and_result98[187]^and_result98[188]^and_result98[189]^and_result98[190]^and_result98[191]^and_result98[192]^and_result98[193]^and_result98[194]^and_result98[195]^and_result98[196]^and_result98[197]^and_result98[198]^and_result98[199]^and_result98[200]^and_result98[201]^and_result98[202]^and_result98[203]^and_result98[204]^and_result98[205]^and_result98[206]^and_result98[207]^and_result98[208]^and_result98[209]^and_result98[210]^and_result98[211]^and_result98[212]^and_result98[213]^and_result98[214]^and_result98[215]^and_result98[216]^and_result98[217]^and_result98[218]^and_result98[219]^and_result98[220]^and_result98[221]^and_result98[222]^and_result98[223]^and_result98[224]^and_result98[225]^and_result98[226]^and_result98[227]^and_result98[228]^and_result98[229]^and_result98[230]^and_result98[231]^and_result98[232]^and_result98[233]^and_result98[234]^and_result98[235]^and_result98[236]^and_result98[237]^and_result98[238]^and_result98[239]^and_result98[240]^and_result98[241]^and_result98[242]^and_result98[243]^and_result98[244]^and_result98[245]^and_result98[246]^and_result98[247]^and_result98[248]^and_result98[249]^and_result98[250]^and_result98[251]^and_result98[252]^and_result98[253]^and_result98[254];
assign key[99]=and_result99[0]^and_result99[1]^and_result99[2]^and_result99[3]^and_result99[4]^and_result99[5]^and_result99[6]^and_result99[7]^and_result99[8]^and_result99[9]^and_result99[10]^and_result99[11]^and_result99[12]^and_result99[13]^and_result99[14]^and_result99[15]^and_result99[16]^and_result99[17]^and_result99[18]^and_result99[19]^and_result99[20]^and_result99[21]^and_result99[22]^and_result99[23]^and_result99[24]^and_result99[25]^and_result99[26]^and_result99[27]^and_result99[28]^and_result99[29]^and_result99[30]^and_result99[31]^and_result99[32]^and_result99[33]^and_result99[34]^and_result99[35]^and_result99[36]^and_result99[37]^and_result99[38]^and_result99[39]^and_result99[40]^and_result99[41]^and_result99[42]^and_result99[43]^and_result99[44]^and_result99[45]^and_result99[46]^and_result99[47]^and_result99[48]^and_result99[49]^and_result99[50]^and_result99[51]^and_result99[52]^and_result99[53]^and_result99[54]^and_result99[55]^and_result99[56]^and_result99[57]^and_result99[58]^and_result99[59]^and_result99[60]^and_result99[61]^and_result99[62]^and_result99[63]^and_result99[64]^and_result99[65]^and_result99[66]^and_result99[67]^and_result99[68]^and_result99[69]^and_result99[70]^and_result99[71]^and_result99[72]^and_result99[73]^and_result99[74]^and_result99[75]^and_result99[76]^and_result99[77]^and_result99[78]^and_result99[79]^and_result99[80]^and_result99[81]^and_result99[82]^and_result99[83]^and_result99[84]^and_result99[85]^and_result99[86]^and_result99[87]^and_result99[88]^and_result99[89]^and_result99[90]^and_result99[91]^and_result99[92]^and_result99[93]^and_result99[94]^and_result99[95]^and_result99[96]^and_result99[97]^and_result99[98]^and_result99[99]^and_result99[100]^and_result99[101]^and_result99[102]^and_result99[103]^and_result99[104]^and_result99[105]^and_result99[106]^and_result99[107]^and_result99[108]^and_result99[109]^and_result99[110]^and_result99[111]^and_result99[112]^and_result99[113]^and_result99[114]^and_result99[115]^and_result99[116]^and_result99[117]^and_result99[118]^and_result99[119]^and_result99[120]^and_result99[121]^and_result99[122]^and_result99[123]^and_result99[124]^and_result99[125]^and_result99[126]^and_result99[127]^and_result99[128]^and_result99[129]^and_result99[130]^and_result99[131]^and_result99[132]^and_result99[133]^and_result99[134]^and_result99[135]^and_result99[136]^and_result99[137]^and_result99[138]^and_result99[139]^and_result99[140]^and_result99[141]^and_result99[142]^and_result99[143]^and_result99[144]^and_result99[145]^and_result99[146]^and_result99[147]^and_result99[148]^and_result99[149]^and_result99[150]^and_result99[151]^and_result99[152]^and_result99[153]^and_result99[154]^and_result99[155]^and_result99[156]^and_result99[157]^and_result99[158]^and_result99[159]^and_result99[160]^and_result99[161]^and_result99[162]^and_result99[163]^and_result99[164]^and_result99[165]^and_result99[166]^and_result99[167]^and_result99[168]^and_result99[169]^and_result99[170]^and_result99[171]^and_result99[172]^and_result99[173]^and_result99[174]^and_result99[175]^and_result99[176]^and_result99[177]^and_result99[178]^and_result99[179]^and_result99[180]^and_result99[181]^and_result99[182]^and_result99[183]^and_result99[184]^and_result99[185]^and_result99[186]^and_result99[187]^and_result99[188]^and_result99[189]^and_result99[190]^and_result99[191]^and_result99[192]^and_result99[193]^and_result99[194]^and_result99[195]^and_result99[196]^and_result99[197]^and_result99[198]^and_result99[199]^and_result99[200]^and_result99[201]^and_result99[202]^and_result99[203]^and_result99[204]^and_result99[205]^and_result99[206]^and_result99[207]^and_result99[208]^and_result99[209]^and_result99[210]^and_result99[211]^and_result99[212]^and_result99[213]^and_result99[214]^and_result99[215]^and_result99[216]^and_result99[217]^and_result99[218]^and_result99[219]^and_result99[220]^and_result99[221]^and_result99[222]^and_result99[223]^and_result99[224]^and_result99[225]^and_result99[226]^and_result99[227]^and_result99[228]^and_result99[229]^and_result99[230]^and_result99[231]^and_result99[232]^and_result99[233]^and_result99[234]^and_result99[235]^and_result99[236]^and_result99[237]^and_result99[238]^and_result99[239]^and_result99[240]^and_result99[241]^and_result99[242]^and_result99[243]^and_result99[244]^and_result99[245]^and_result99[246]^and_result99[247]^and_result99[248]^and_result99[249]^and_result99[250]^and_result99[251]^and_result99[252]^and_result99[253]^and_result99[254];
assign key[100]=and_result100[0]^and_result100[1]^and_result100[2]^and_result100[3]^and_result100[4]^and_result100[5]^and_result100[6]^and_result100[7]^and_result100[8]^and_result100[9]^and_result100[10]^and_result100[11]^and_result100[12]^and_result100[13]^and_result100[14]^and_result100[15]^and_result100[16]^and_result100[17]^and_result100[18]^and_result100[19]^and_result100[20]^and_result100[21]^and_result100[22]^and_result100[23]^and_result100[24]^and_result100[25]^and_result100[26]^and_result100[27]^and_result100[28]^and_result100[29]^and_result100[30]^and_result100[31]^and_result100[32]^and_result100[33]^and_result100[34]^and_result100[35]^and_result100[36]^and_result100[37]^and_result100[38]^and_result100[39]^and_result100[40]^and_result100[41]^and_result100[42]^and_result100[43]^and_result100[44]^and_result100[45]^and_result100[46]^and_result100[47]^and_result100[48]^and_result100[49]^and_result100[50]^and_result100[51]^and_result100[52]^and_result100[53]^and_result100[54]^and_result100[55]^and_result100[56]^and_result100[57]^and_result100[58]^and_result100[59]^and_result100[60]^and_result100[61]^and_result100[62]^and_result100[63]^and_result100[64]^and_result100[65]^and_result100[66]^and_result100[67]^and_result100[68]^and_result100[69]^and_result100[70]^and_result100[71]^and_result100[72]^and_result100[73]^and_result100[74]^and_result100[75]^and_result100[76]^and_result100[77]^and_result100[78]^and_result100[79]^and_result100[80]^and_result100[81]^and_result100[82]^and_result100[83]^and_result100[84]^and_result100[85]^and_result100[86]^and_result100[87]^and_result100[88]^and_result100[89]^and_result100[90]^and_result100[91]^and_result100[92]^and_result100[93]^and_result100[94]^and_result100[95]^and_result100[96]^and_result100[97]^and_result100[98]^and_result100[99]^and_result100[100]^and_result100[101]^and_result100[102]^and_result100[103]^and_result100[104]^and_result100[105]^and_result100[106]^and_result100[107]^and_result100[108]^and_result100[109]^and_result100[110]^and_result100[111]^and_result100[112]^and_result100[113]^and_result100[114]^and_result100[115]^and_result100[116]^and_result100[117]^and_result100[118]^and_result100[119]^and_result100[120]^and_result100[121]^and_result100[122]^and_result100[123]^and_result100[124]^and_result100[125]^and_result100[126]^and_result100[127]^and_result100[128]^and_result100[129]^and_result100[130]^and_result100[131]^and_result100[132]^and_result100[133]^and_result100[134]^and_result100[135]^and_result100[136]^and_result100[137]^and_result100[138]^and_result100[139]^and_result100[140]^and_result100[141]^and_result100[142]^and_result100[143]^and_result100[144]^and_result100[145]^and_result100[146]^and_result100[147]^and_result100[148]^and_result100[149]^and_result100[150]^and_result100[151]^and_result100[152]^and_result100[153]^and_result100[154]^and_result100[155]^and_result100[156]^and_result100[157]^and_result100[158]^and_result100[159]^and_result100[160]^and_result100[161]^and_result100[162]^and_result100[163]^and_result100[164]^and_result100[165]^and_result100[166]^and_result100[167]^and_result100[168]^and_result100[169]^and_result100[170]^and_result100[171]^and_result100[172]^and_result100[173]^and_result100[174]^and_result100[175]^and_result100[176]^and_result100[177]^and_result100[178]^and_result100[179]^and_result100[180]^and_result100[181]^and_result100[182]^and_result100[183]^and_result100[184]^and_result100[185]^and_result100[186]^and_result100[187]^and_result100[188]^and_result100[189]^and_result100[190]^and_result100[191]^and_result100[192]^and_result100[193]^and_result100[194]^and_result100[195]^and_result100[196]^and_result100[197]^and_result100[198]^and_result100[199]^and_result100[200]^and_result100[201]^and_result100[202]^and_result100[203]^and_result100[204]^and_result100[205]^and_result100[206]^and_result100[207]^and_result100[208]^and_result100[209]^and_result100[210]^and_result100[211]^and_result100[212]^and_result100[213]^and_result100[214]^and_result100[215]^and_result100[216]^and_result100[217]^and_result100[218]^and_result100[219]^and_result100[220]^and_result100[221]^and_result100[222]^and_result100[223]^and_result100[224]^and_result100[225]^and_result100[226]^and_result100[227]^and_result100[228]^and_result100[229]^and_result100[230]^and_result100[231]^and_result100[232]^and_result100[233]^and_result100[234]^and_result100[235]^and_result100[236]^and_result100[237]^and_result100[238]^and_result100[239]^and_result100[240]^and_result100[241]^and_result100[242]^and_result100[243]^and_result100[244]^and_result100[245]^and_result100[246]^and_result100[247]^and_result100[248]^and_result100[249]^and_result100[250]^and_result100[251]^and_result100[252]^and_result100[253]^and_result100[254];
assign key[101]=and_result101[0]^and_result101[1]^and_result101[2]^and_result101[3]^and_result101[4]^and_result101[5]^and_result101[6]^and_result101[7]^and_result101[8]^and_result101[9]^and_result101[10]^and_result101[11]^and_result101[12]^and_result101[13]^and_result101[14]^and_result101[15]^and_result101[16]^and_result101[17]^and_result101[18]^and_result101[19]^and_result101[20]^and_result101[21]^and_result101[22]^and_result101[23]^and_result101[24]^and_result101[25]^and_result101[26]^and_result101[27]^and_result101[28]^and_result101[29]^and_result101[30]^and_result101[31]^and_result101[32]^and_result101[33]^and_result101[34]^and_result101[35]^and_result101[36]^and_result101[37]^and_result101[38]^and_result101[39]^and_result101[40]^and_result101[41]^and_result101[42]^and_result101[43]^and_result101[44]^and_result101[45]^and_result101[46]^and_result101[47]^and_result101[48]^and_result101[49]^and_result101[50]^and_result101[51]^and_result101[52]^and_result101[53]^and_result101[54]^and_result101[55]^and_result101[56]^and_result101[57]^and_result101[58]^and_result101[59]^and_result101[60]^and_result101[61]^and_result101[62]^and_result101[63]^and_result101[64]^and_result101[65]^and_result101[66]^and_result101[67]^and_result101[68]^and_result101[69]^and_result101[70]^and_result101[71]^and_result101[72]^and_result101[73]^and_result101[74]^and_result101[75]^and_result101[76]^and_result101[77]^and_result101[78]^and_result101[79]^and_result101[80]^and_result101[81]^and_result101[82]^and_result101[83]^and_result101[84]^and_result101[85]^and_result101[86]^and_result101[87]^and_result101[88]^and_result101[89]^and_result101[90]^and_result101[91]^and_result101[92]^and_result101[93]^and_result101[94]^and_result101[95]^and_result101[96]^and_result101[97]^and_result101[98]^and_result101[99]^and_result101[100]^and_result101[101]^and_result101[102]^and_result101[103]^and_result101[104]^and_result101[105]^and_result101[106]^and_result101[107]^and_result101[108]^and_result101[109]^and_result101[110]^and_result101[111]^and_result101[112]^and_result101[113]^and_result101[114]^and_result101[115]^and_result101[116]^and_result101[117]^and_result101[118]^and_result101[119]^and_result101[120]^and_result101[121]^and_result101[122]^and_result101[123]^and_result101[124]^and_result101[125]^and_result101[126]^and_result101[127]^and_result101[128]^and_result101[129]^and_result101[130]^and_result101[131]^and_result101[132]^and_result101[133]^and_result101[134]^and_result101[135]^and_result101[136]^and_result101[137]^and_result101[138]^and_result101[139]^and_result101[140]^and_result101[141]^and_result101[142]^and_result101[143]^and_result101[144]^and_result101[145]^and_result101[146]^and_result101[147]^and_result101[148]^and_result101[149]^and_result101[150]^and_result101[151]^and_result101[152]^and_result101[153]^and_result101[154]^and_result101[155]^and_result101[156]^and_result101[157]^and_result101[158]^and_result101[159]^and_result101[160]^and_result101[161]^and_result101[162]^and_result101[163]^and_result101[164]^and_result101[165]^and_result101[166]^and_result101[167]^and_result101[168]^and_result101[169]^and_result101[170]^and_result101[171]^and_result101[172]^and_result101[173]^and_result101[174]^and_result101[175]^and_result101[176]^and_result101[177]^and_result101[178]^and_result101[179]^and_result101[180]^and_result101[181]^and_result101[182]^and_result101[183]^and_result101[184]^and_result101[185]^and_result101[186]^and_result101[187]^and_result101[188]^and_result101[189]^and_result101[190]^and_result101[191]^and_result101[192]^and_result101[193]^and_result101[194]^and_result101[195]^and_result101[196]^and_result101[197]^and_result101[198]^and_result101[199]^and_result101[200]^and_result101[201]^and_result101[202]^and_result101[203]^and_result101[204]^and_result101[205]^and_result101[206]^and_result101[207]^and_result101[208]^and_result101[209]^and_result101[210]^and_result101[211]^and_result101[212]^and_result101[213]^and_result101[214]^and_result101[215]^and_result101[216]^and_result101[217]^and_result101[218]^and_result101[219]^and_result101[220]^and_result101[221]^and_result101[222]^and_result101[223]^and_result101[224]^and_result101[225]^and_result101[226]^and_result101[227]^and_result101[228]^and_result101[229]^and_result101[230]^and_result101[231]^and_result101[232]^and_result101[233]^and_result101[234]^and_result101[235]^and_result101[236]^and_result101[237]^and_result101[238]^and_result101[239]^and_result101[240]^and_result101[241]^and_result101[242]^and_result101[243]^and_result101[244]^and_result101[245]^and_result101[246]^and_result101[247]^and_result101[248]^and_result101[249]^and_result101[250]^and_result101[251]^and_result101[252]^and_result101[253]^and_result101[254];
assign key[102]=and_result102[0]^and_result102[1]^and_result102[2]^and_result102[3]^and_result102[4]^and_result102[5]^and_result102[6]^and_result102[7]^and_result102[8]^and_result102[9]^and_result102[10]^and_result102[11]^and_result102[12]^and_result102[13]^and_result102[14]^and_result102[15]^and_result102[16]^and_result102[17]^and_result102[18]^and_result102[19]^and_result102[20]^and_result102[21]^and_result102[22]^and_result102[23]^and_result102[24]^and_result102[25]^and_result102[26]^and_result102[27]^and_result102[28]^and_result102[29]^and_result102[30]^and_result102[31]^and_result102[32]^and_result102[33]^and_result102[34]^and_result102[35]^and_result102[36]^and_result102[37]^and_result102[38]^and_result102[39]^and_result102[40]^and_result102[41]^and_result102[42]^and_result102[43]^and_result102[44]^and_result102[45]^and_result102[46]^and_result102[47]^and_result102[48]^and_result102[49]^and_result102[50]^and_result102[51]^and_result102[52]^and_result102[53]^and_result102[54]^and_result102[55]^and_result102[56]^and_result102[57]^and_result102[58]^and_result102[59]^and_result102[60]^and_result102[61]^and_result102[62]^and_result102[63]^and_result102[64]^and_result102[65]^and_result102[66]^and_result102[67]^and_result102[68]^and_result102[69]^and_result102[70]^and_result102[71]^and_result102[72]^and_result102[73]^and_result102[74]^and_result102[75]^and_result102[76]^and_result102[77]^and_result102[78]^and_result102[79]^and_result102[80]^and_result102[81]^and_result102[82]^and_result102[83]^and_result102[84]^and_result102[85]^and_result102[86]^and_result102[87]^and_result102[88]^and_result102[89]^and_result102[90]^and_result102[91]^and_result102[92]^and_result102[93]^and_result102[94]^and_result102[95]^and_result102[96]^and_result102[97]^and_result102[98]^and_result102[99]^and_result102[100]^and_result102[101]^and_result102[102]^and_result102[103]^and_result102[104]^and_result102[105]^and_result102[106]^and_result102[107]^and_result102[108]^and_result102[109]^and_result102[110]^and_result102[111]^and_result102[112]^and_result102[113]^and_result102[114]^and_result102[115]^and_result102[116]^and_result102[117]^and_result102[118]^and_result102[119]^and_result102[120]^and_result102[121]^and_result102[122]^and_result102[123]^and_result102[124]^and_result102[125]^and_result102[126]^and_result102[127]^and_result102[128]^and_result102[129]^and_result102[130]^and_result102[131]^and_result102[132]^and_result102[133]^and_result102[134]^and_result102[135]^and_result102[136]^and_result102[137]^and_result102[138]^and_result102[139]^and_result102[140]^and_result102[141]^and_result102[142]^and_result102[143]^and_result102[144]^and_result102[145]^and_result102[146]^and_result102[147]^and_result102[148]^and_result102[149]^and_result102[150]^and_result102[151]^and_result102[152]^and_result102[153]^and_result102[154]^and_result102[155]^and_result102[156]^and_result102[157]^and_result102[158]^and_result102[159]^and_result102[160]^and_result102[161]^and_result102[162]^and_result102[163]^and_result102[164]^and_result102[165]^and_result102[166]^and_result102[167]^and_result102[168]^and_result102[169]^and_result102[170]^and_result102[171]^and_result102[172]^and_result102[173]^and_result102[174]^and_result102[175]^and_result102[176]^and_result102[177]^and_result102[178]^and_result102[179]^and_result102[180]^and_result102[181]^and_result102[182]^and_result102[183]^and_result102[184]^and_result102[185]^and_result102[186]^and_result102[187]^and_result102[188]^and_result102[189]^and_result102[190]^and_result102[191]^and_result102[192]^and_result102[193]^and_result102[194]^and_result102[195]^and_result102[196]^and_result102[197]^and_result102[198]^and_result102[199]^and_result102[200]^and_result102[201]^and_result102[202]^and_result102[203]^and_result102[204]^and_result102[205]^and_result102[206]^and_result102[207]^and_result102[208]^and_result102[209]^and_result102[210]^and_result102[211]^and_result102[212]^and_result102[213]^and_result102[214]^and_result102[215]^and_result102[216]^and_result102[217]^and_result102[218]^and_result102[219]^and_result102[220]^and_result102[221]^and_result102[222]^and_result102[223]^and_result102[224]^and_result102[225]^and_result102[226]^and_result102[227]^and_result102[228]^and_result102[229]^and_result102[230]^and_result102[231]^and_result102[232]^and_result102[233]^and_result102[234]^and_result102[235]^and_result102[236]^and_result102[237]^and_result102[238]^and_result102[239]^and_result102[240]^and_result102[241]^and_result102[242]^and_result102[243]^and_result102[244]^and_result102[245]^and_result102[246]^and_result102[247]^and_result102[248]^and_result102[249]^and_result102[250]^and_result102[251]^and_result102[252]^and_result102[253]^and_result102[254];
assign key[103]=and_result103[0]^and_result103[1]^and_result103[2]^and_result103[3]^and_result103[4]^and_result103[5]^and_result103[6]^and_result103[7]^and_result103[8]^and_result103[9]^and_result103[10]^and_result103[11]^and_result103[12]^and_result103[13]^and_result103[14]^and_result103[15]^and_result103[16]^and_result103[17]^and_result103[18]^and_result103[19]^and_result103[20]^and_result103[21]^and_result103[22]^and_result103[23]^and_result103[24]^and_result103[25]^and_result103[26]^and_result103[27]^and_result103[28]^and_result103[29]^and_result103[30]^and_result103[31]^and_result103[32]^and_result103[33]^and_result103[34]^and_result103[35]^and_result103[36]^and_result103[37]^and_result103[38]^and_result103[39]^and_result103[40]^and_result103[41]^and_result103[42]^and_result103[43]^and_result103[44]^and_result103[45]^and_result103[46]^and_result103[47]^and_result103[48]^and_result103[49]^and_result103[50]^and_result103[51]^and_result103[52]^and_result103[53]^and_result103[54]^and_result103[55]^and_result103[56]^and_result103[57]^and_result103[58]^and_result103[59]^and_result103[60]^and_result103[61]^and_result103[62]^and_result103[63]^and_result103[64]^and_result103[65]^and_result103[66]^and_result103[67]^and_result103[68]^and_result103[69]^and_result103[70]^and_result103[71]^and_result103[72]^and_result103[73]^and_result103[74]^and_result103[75]^and_result103[76]^and_result103[77]^and_result103[78]^and_result103[79]^and_result103[80]^and_result103[81]^and_result103[82]^and_result103[83]^and_result103[84]^and_result103[85]^and_result103[86]^and_result103[87]^and_result103[88]^and_result103[89]^and_result103[90]^and_result103[91]^and_result103[92]^and_result103[93]^and_result103[94]^and_result103[95]^and_result103[96]^and_result103[97]^and_result103[98]^and_result103[99]^and_result103[100]^and_result103[101]^and_result103[102]^and_result103[103]^and_result103[104]^and_result103[105]^and_result103[106]^and_result103[107]^and_result103[108]^and_result103[109]^and_result103[110]^and_result103[111]^and_result103[112]^and_result103[113]^and_result103[114]^and_result103[115]^and_result103[116]^and_result103[117]^and_result103[118]^and_result103[119]^and_result103[120]^and_result103[121]^and_result103[122]^and_result103[123]^and_result103[124]^and_result103[125]^and_result103[126]^and_result103[127]^and_result103[128]^and_result103[129]^and_result103[130]^and_result103[131]^and_result103[132]^and_result103[133]^and_result103[134]^and_result103[135]^and_result103[136]^and_result103[137]^and_result103[138]^and_result103[139]^and_result103[140]^and_result103[141]^and_result103[142]^and_result103[143]^and_result103[144]^and_result103[145]^and_result103[146]^and_result103[147]^and_result103[148]^and_result103[149]^and_result103[150]^and_result103[151]^and_result103[152]^and_result103[153]^and_result103[154]^and_result103[155]^and_result103[156]^and_result103[157]^and_result103[158]^and_result103[159]^and_result103[160]^and_result103[161]^and_result103[162]^and_result103[163]^and_result103[164]^and_result103[165]^and_result103[166]^and_result103[167]^and_result103[168]^and_result103[169]^and_result103[170]^and_result103[171]^and_result103[172]^and_result103[173]^and_result103[174]^and_result103[175]^and_result103[176]^and_result103[177]^and_result103[178]^and_result103[179]^and_result103[180]^and_result103[181]^and_result103[182]^and_result103[183]^and_result103[184]^and_result103[185]^and_result103[186]^and_result103[187]^and_result103[188]^and_result103[189]^and_result103[190]^and_result103[191]^and_result103[192]^and_result103[193]^and_result103[194]^and_result103[195]^and_result103[196]^and_result103[197]^and_result103[198]^and_result103[199]^and_result103[200]^and_result103[201]^and_result103[202]^and_result103[203]^and_result103[204]^and_result103[205]^and_result103[206]^and_result103[207]^and_result103[208]^and_result103[209]^and_result103[210]^and_result103[211]^and_result103[212]^and_result103[213]^and_result103[214]^and_result103[215]^and_result103[216]^and_result103[217]^and_result103[218]^and_result103[219]^and_result103[220]^and_result103[221]^and_result103[222]^and_result103[223]^and_result103[224]^and_result103[225]^and_result103[226]^and_result103[227]^and_result103[228]^and_result103[229]^and_result103[230]^and_result103[231]^and_result103[232]^and_result103[233]^and_result103[234]^and_result103[235]^and_result103[236]^and_result103[237]^and_result103[238]^and_result103[239]^and_result103[240]^and_result103[241]^and_result103[242]^and_result103[243]^and_result103[244]^and_result103[245]^and_result103[246]^and_result103[247]^and_result103[248]^and_result103[249]^and_result103[250]^and_result103[251]^and_result103[252]^and_result103[253]^and_result103[254];
assign key[104]=and_result104[0]^and_result104[1]^and_result104[2]^and_result104[3]^and_result104[4]^and_result104[5]^and_result104[6]^and_result104[7]^and_result104[8]^and_result104[9]^and_result104[10]^and_result104[11]^and_result104[12]^and_result104[13]^and_result104[14]^and_result104[15]^and_result104[16]^and_result104[17]^and_result104[18]^and_result104[19]^and_result104[20]^and_result104[21]^and_result104[22]^and_result104[23]^and_result104[24]^and_result104[25]^and_result104[26]^and_result104[27]^and_result104[28]^and_result104[29]^and_result104[30]^and_result104[31]^and_result104[32]^and_result104[33]^and_result104[34]^and_result104[35]^and_result104[36]^and_result104[37]^and_result104[38]^and_result104[39]^and_result104[40]^and_result104[41]^and_result104[42]^and_result104[43]^and_result104[44]^and_result104[45]^and_result104[46]^and_result104[47]^and_result104[48]^and_result104[49]^and_result104[50]^and_result104[51]^and_result104[52]^and_result104[53]^and_result104[54]^and_result104[55]^and_result104[56]^and_result104[57]^and_result104[58]^and_result104[59]^and_result104[60]^and_result104[61]^and_result104[62]^and_result104[63]^and_result104[64]^and_result104[65]^and_result104[66]^and_result104[67]^and_result104[68]^and_result104[69]^and_result104[70]^and_result104[71]^and_result104[72]^and_result104[73]^and_result104[74]^and_result104[75]^and_result104[76]^and_result104[77]^and_result104[78]^and_result104[79]^and_result104[80]^and_result104[81]^and_result104[82]^and_result104[83]^and_result104[84]^and_result104[85]^and_result104[86]^and_result104[87]^and_result104[88]^and_result104[89]^and_result104[90]^and_result104[91]^and_result104[92]^and_result104[93]^and_result104[94]^and_result104[95]^and_result104[96]^and_result104[97]^and_result104[98]^and_result104[99]^and_result104[100]^and_result104[101]^and_result104[102]^and_result104[103]^and_result104[104]^and_result104[105]^and_result104[106]^and_result104[107]^and_result104[108]^and_result104[109]^and_result104[110]^and_result104[111]^and_result104[112]^and_result104[113]^and_result104[114]^and_result104[115]^and_result104[116]^and_result104[117]^and_result104[118]^and_result104[119]^and_result104[120]^and_result104[121]^and_result104[122]^and_result104[123]^and_result104[124]^and_result104[125]^and_result104[126]^and_result104[127]^and_result104[128]^and_result104[129]^and_result104[130]^and_result104[131]^and_result104[132]^and_result104[133]^and_result104[134]^and_result104[135]^and_result104[136]^and_result104[137]^and_result104[138]^and_result104[139]^and_result104[140]^and_result104[141]^and_result104[142]^and_result104[143]^and_result104[144]^and_result104[145]^and_result104[146]^and_result104[147]^and_result104[148]^and_result104[149]^and_result104[150]^and_result104[151]^and_result104[152]^and_result104[153]^and_result104[154]^and_result104[155]^and_result104[156]^and_result104[157]^and_result104[158]^and_result104[159]^and_result104[160]^and_result104[161]^and_result104[162]^and_result104[163]^and_result104[164]^and_result104[165]^and_result104[166]^and_result104[167]^and_result104[168]^and_result104[169]^and_result104[170]^and_result104[171]^and_result104[172]^and_result104[173]^and_result104[174]^and_result104[175]^and_result104[176]^and_result104[177]^and_result104[178]^and_result104[179]^and_result104[180]^and_result104[181]^and_result104[182]^and_result104[183]^and_result104[184]^and_result104[185]^and_result104[186]^and_result104[187]^and_result104[188]^and_result104[189]^and_result104[190]^and_result104[191]^and_result104[192]^and_result104[193]^and_result104[194]^and_result104[195]^and_result104[196]^and_result104[197]^and_result104[198]^and_result104[199]^and_result104[200]^and_result104[201]^and_result104[202]^and_result104[203]^and_result104[204]^and_result104[205]^and_result104[206]^and_result104[207]^and_result104[208]^and_result104[209]^and_result104[210]^and_result104[211]^and_result104[212]^and_result104[213]^and_result104[214]^and_result104[215]^and_result104[216]^and_result104[217]^and_result104[218]^and_result104[219]^and_result104[220]^and_result104[221]^and_result104[222]^and_result104[223]^and_result104[224]^and_result104[225]^and_result104[226]^and_result104[227]^and_result104[228]^and_result104[229]^and_result104[230]^and_result104[231]^and_result104[232]^and_result104[233]^and_result104[234]^and_result104[235]^and_result104[236]^and_result104[237]^and_result104[238]^and_result104[239]^and_result104[240]^and_result104[241]^and_result104[242]^and_result104[243]^and_result104[244]^and_result104[245]^and_result104[246]^and_result104[247]^and_result104[248]^and_result104[249]^and_result104[250]^and_result104[251]^and_result104[252]^and_result104[253]^and_result104[254];
assign key[105]=and_result105[0]^and_result105[1]^and_result105[2]^and_result105[3]^and_result105[4]^and_result105[5]^and_result105[6]^and_result105[7]^and_result105[8]^and_result105[9]^and_result105[10]^and_result105[11]^and_result105[12]^and_result105[13]^and_result105[14]^and_result105[15]^and_result105[16]^and_result105[17]^and_result105[18]^and_result105[19]^and_result105[20]^and_result105[21]^and_result105[22]^and_result105[23]^and_result105[24]^and_result105[25]^and_result105[26]^and_result105[27]^and_result105[28]^and_result105[29]^and_result105[30]^and_result105[31]^and_result105[32]^and_result105[33]^and_result105[34]^and_result105[35]^and_result105[36]^and_result105[37]^and_result105[38]^and_result105[39]^and_result105[40]^and_result105[41]^and_result105[42]^and_result105[43]^and_result105[44]^and_result105[45]^and_result105[46]^and_result105[47]^and_result105[48]^and_result105[49]^and_result105[50]^and_result105[51]^and_result105[52]^and_result105[53]^and_result105[54]^and_result105[55]^and_result105[56]^and_result105[57]^and_result105[58]^and_result105[59]^and_result105[60]^and_result105[61]^and_result105[62]^and_result105[63]^and_result105[64]^and_result105[65]^and_result105[66]^and_result105[67]^and_result105[68]^and_result105[69]^and_result105[70]^and_result105[71]^and_result105[72]^and_result105[73]^and_result105[74]^and_result105[75]^and_result105[76]^and_result105[77]^and_result105[78]^and_result105[79]^and_result105[80]^and_result105[81]^and_result105[82]^and_result105[83]^and_result105[84]^and_result105[85]^and_result105[86]^and_result105[87]^and_result105[88]^and_result105[89]^and_result105[90]^and_result105[91]^and_result105[92]^and_result105[93]^and_result105[94]^and_result105[95]^and_result105[96]^and_result105[97]^and_result105[98]^and_result105[99]^and_result105[100]^and_result105[101]^and_result105[102]^and_result105[103]^and_result105[104]^and_result105[105]^and_result105[106]^and_result105[107]^and_result105[108]^and_result105[109]^and_result105[110]^and_result105[111]^and_result105[112]^and_result105[113]^and_result105[114]^and_result105[115]^and_result105[116]^and_result105[117]^and_result105[118]^and_result105[119]^and_result105[120]^and_result105[121]^and_result105[122]^and_result105[123]^and_result105[124]^and_result105[125]^and_result105[126]^and_result105[127]^and_result105[128]^and_result105[129]^and_result105[130]^and_result105[131]^and_result105[132]^and_result105[133]^and_result105[134]^and_result105[135]^and_result105[136]^and_result105[137]^and_result105[138]^and_result105[139]^and_result105[140]^and_result105[141]^and_result105[142]^and_result105[143]^and_result105[144]^and_result105[145]^and_result105[146]^and_result105[147]^and_result105[148]^and_result105[149]^and_result105[150]^and_result105[151]^and_result105[152]^and_result105[153]^and_result105[154]^and_result105[155]^and_result105[156]^and_result105[157]^and_result105[158]^and_result105[159]^and_result105[160]^and_result105[161]^and_result105[162]^and_result105[163]^and_result105[164]^and_result105[165]^and_result105[166]^and_result105[167]^and_result105[168]^and_result105[169]^and_result105[170]^and_result105[171]^and_result105[172]^and_result105[173]^and_result105[174]^and_result105[175]^and_result105[176]^and_result105[177]^and_result105[178]^and_result105[179]^and_result105[180]^and_result105[181]^and_result105[182]^and_result105[183]^and_result105[184]^and_result105[185]^and_result105[186]^and_result105[187]^and_result105[188]^and_result105[189]^and_result105[190]^and_result105[191]^and_result105[192]^and_result105[193]^and_result105[194]^and_result105[195]^and_result105[196]^and_result105[197]^and_result105[198]^and_result105[199]^and_result105[200]^and_result105[201]^and_result105[202]^and_result105[203]^and_result105[204]^and_result105[205]^and_result105[206]^and_result105[207]^and_result105[208]^and_result105[209]^and_result105[210]^and_result105[211]^and_result105[212]^and_result105[213]^and_result105[214]^and_result105[215]^and_result105[216]^and_result105[217]^and_result105[218]^and_result105[219]^and_result105[220]^and_result105[221]^and_result105[222]^and_result105[223]^and_result105[224]^and_result105[225]^and_result105[226]^and_result105[227]^and_result105[228]^and_result105[229]^and_result105[230]^and_result105[231]^and_result105[232]^and_result105[233]^and_result105[234]^and_result105[235]^and_result105[236]^and_result105[237]^and_result105[238]^and_result105[239]^and_result105[240]^and_result105[241]^and_result105[242]^and_result105[243]^and_result105[244]^and_result105[245]^and_result105[246]^and_result105[247]^and_result105[248]^and_result105[249]^and_result105[250]^and_result105[251]^and_result105[252]^and_result105[253]^and_result105[254];
assign key[106]=and_result106[0]^and_result106[1]^and_result106[2]^and_result106[3]^and_result106[4]^and_result106[5]^and_result106[6]^and_result106[7]^and_result106[8]^and_result106[9]^and_result106[10]^and_result106[11]^and_result106[12]^and_result106[13]^and_result106[14]^and_result106[15]^and_result106[16]^and_result106[17]^and_result106[18]^and_result106[19]^and_result106[20]^and_result106[21]^and_result106[22]^and_result106[23]^and_result106[24]^and_result106[25]^and_result106[26]^and_result106[27]^and_result106[28]^and_result106[29]^and_result106[30]^and_result106[31]^and_result106[32]^and_result106[33]^and_result106[34]^and_result106[35]^and_result106[36]^and_result106[37]^and_result106[38]^and_result106[39]^and_result106[40]^and_result106[41]^and_result106[42]^and_result106[43]^and_result106[44]^and_result106[45]^and_result106[46]^and_result106[47]^and_result106[48]^and_result106[49]^and_result106[50]^and_result106[51]^and_result106[52]^and_result106[53]^and_result106[54]^and_result106[55]^and_result106[56]^and_result106[57]^and_result106[58]^and_result106[59]^and_result106[60]^and_result106[61]^and_result106[62]^and_result106[63]^and_result106[64]^and_result106[65]^and_result106[66]^and_result106[67]^and_result106[68]^and_result106[69]^and_result106[70]^and_result106[71]^and_result106[72]^and_result106[73]^and_result106[74]^and_result106[75]^and_result106[76]^and_result106[77]^and_result106[78]^and_result106[79]^and_result106[80]^and_result106[81]^and_result106[82]^and_result106[83]^and_result106[84]^and_result106[85]^and_result106[86]^and_result106[87]^and_result106[88]^and_result106[89]^and_result106[90]^and_result106[91]^and_result106[92]^and_result106[93]^and_result106[94]^and_result106[95]^and_result106[96]^and_result106[97]^and_result106[98]^and_result106[99]^and_result106[100]^and_result106[101]^and_result106[102]^and_result106[103]^and_result106[104]^and_result106[105]^and_result106[106]^and_result106[107]^and_result106[108]^and_result106[109]^and_result106[110]^and_result106[111]^and_result106[112]^and_result106[113]^and_result106[114]^and_result106[115]^and_result106[116]^and_result106[117]^and_result106[118]^and_result106[119]^and_result106[120]^and_result106[121]^and_result106[122]^and_result106[123]^and_result106[124]^and_result106[125]^and_result106[126]^and_result106[127]^and_result106[128]^and_result106[129]^and_result106[130]^and_result106[131]^and_result106[132]^and_result106[133]^and_result106[134]^and_result106[135]^and_result106[136]^and_result106[137]^and_result106[138]^and_result106[139]^and_result106[140]^and_result106[141]^and_result106[142]^and_result106[143]^and_result106[144]^and_result106[145]^and_result106[146]^and_result106[147]^and_result106[148]^and_result106[149]^and_result106[150]^and_result106[151]^and_result106[152]^and_result106[153]^and_result106[154]^and_result106[155]^and_result106[156]^and_result106[157]^and_result106[158]^and_result106[159]^and_result106[160]^and_result106[161]^and_result106[162]^and_result106[163]^and_result106[164]^and_result106[165]^and_result106[166]^and_result106[167]^and_result106[168]^and_result106[169]^and_result106[170]^and_result106[171]^and_result106[172]^and_result106[173]^and_result106[174]^and_result106[175]^and_result106[176]^and_result106[177]^and_result106[178]^and_result106[179]^and_result106[180]^and_result106[181]^and_result106[182]^and_result106[183]^and_result106[184]^and_result106[185]^and_result106[186]^and_result106[187]^and_result106[188]^and_result106[189]^and_result106[190]^and_result106[191]^and_result106[192]^and_result106[193]^and_result106[194]^and_result106[195]^and_result106[196]^and_result106[197]^and_result106[198]^and_result106[199]^and_result106[200]^and_result106[201]^and_result106[202]^and_result106[203]^and_result106[204]^and_result106[205]^and_result106[206]^and_result106[207]^and_result106[208]^and_result106[209]^and_result106[210]^and_result106[211]^and_result106[212]^and_result106[213]^and_result106[214]^and_result106[215]^and_result106[216]^and_result106[217]^and_result106[218]^and_result106[219]^and_result106[220]^and_result106[221]^and_result106[222]^and_result106[223]^and_result106[224]^and_result106[225]^and_result106[226]^and_result106[227]^and_result106[228]^and_result106[229]^and_result106[230]^and_result106[231]^and_result106[232]^and_result106[233]^and_result106[234]^and_result106[235]^and_result106[236]^and_result106[237]^and_result106[238]^and_result106[239]^and_result106[240]^and_result106[241]^and_result106[242]^and_result106[243]^and_result106[244]^and_result106[245]^and_result106[246]^and_result106[247]^and_result106[248]^and_result106[249]^and_result106[250]^and_result106[251]^and_result106[252]^and_result106[253]^and_result106[254];
assign key[107]=and_result107[0]^and_result107[1]^and_result107[2]^and_result107[3]^and_result107[4]^and_result107[5]^and_result107[6]^and_result107[7]^and_result107[8]^and_result107[9]^and_result107[10]^and_result107[11]^and_result107[12]^and_result107[13]^and_result107[14]^and_result107[15]^and_result107[16]^and_result107[17]^and_result107[18]^and_result107[19]^and_result107[20]^and_result107[21]^and_result107[22]^and_result107[23]^and_result107[24]^and_result107[25]^and_result107[26]^and_result107[27]^and_result107[28]^and_result107[29]^and_result107[30]^and_result107[31]^and_result107[32]^and_result107[33]^and_result107[34]^and_result107[35]^and_result107[36]^and_result107[37]^and_result107[38]^and_result107[39]^and_result107[40]^and_result107[41]^and_result107[42]^and_result107[43]^and_result107[44]^and_result107[45]^and_result107[46]^and_result107[47]^and_result107[48]^and_result107[49]^and_result107[50]^and_result107[51]^and_result107[52]^and_result107[53]^and_result107[54]^and_result107[55]^and_result107[56]^and_result107[57]^and_result107[58]^and_result107[59]^and_result107[60]^and_result107[61]^and_result107[62]^and_result107[63]^and_result107[64]^and_result107[65]^and_result107[66]^and_result107[67]^and_result107[68]^and_result107[69]^and_result107[70]^and_result107[71]^and_result107[72]^and_result107[73]^and_result107[74]^and_result107[75]^and_result107[76]^and_result107[77]^and_result107[78]^and_result107[79]^and_result107[80]^and_result107[81]^and_result107[82]^and_result107[83]^and_result107[84]^and_result107[85]^and_result107[86]^and_result107[87]^and_result107[88]^and_result107[89]^and_result107[90]^and_result107[91]^and_result107[92]^and_result107[93]^and_result107[94]^and_result107[95]^and_result107[96]^and_result107[97]^and_result107[98]^and_result107[99]^and_result107[100]^and_result107[101]^and_result107[102]^and_result107[103]^and_result107[104]^and_result107[105]^and_result107[106]^and_result107[107]^and_result107[108]^and_result107[109]^and_result107[110]^and_result107[111]^and_result107[112]^and_result107[113]^and_result107[114]^and_result107[115]^and_result107[116]^and_result107[117]^and_result107[118]^and_result107[119]^and_result107[120]^and_result107[121]^and_result107[122]^and_result107[123]^and_result107[124]^and_result107[125]^and_result107[126]^and_result107[127]^and_result107[128]^and_result107[129]^and_result107[130]^and_result107[131]^and_result107[132]^and_result107[133]^and_result107[134]^and_result107[135]^and_result107[136]^and_result107[137]^and_result107[138]^and_result107[139]^and_result107[140]^and_result107[141]^and_result107[142]^and_result107[143]^and_result107[144]^and_result107[145]^and_result107[146]^and_result107[147]^and_result107[148]^and_result107[149]^and_result107[150]^and_result107[151]^and_result107[152]^and_result107[153]^and_result107[154]^and_result107[155]^and_result107[156]^and_result107[157]^and_result107[158]^and_result107[159]^and_result107[160]^and_result107[161]^and_result107[162]^and_result107[163]^and_result107[164]^and_result107[165]^and_result107[166]^and_result107[167]^and_result107[168]^and_result107[169]^and_result107[170]^and_result107[171]^and_result107[172]^and_result107[173]^and_result107[174]^and_result107[175]^and_result107[176]^and_result107[177]^and_result107[178]^and_result107[179]^and_result107[180]^and_result107[181]^and_result107[182]^and_result107[183]^and_result107[184]^and_result107[185]^and_result107[186]^and_result107[187]^and_result107[188]^and_result107[189]^and_result107[190]^and_result107[191]^and_result107[192]^and_result107[193]^and_result107[194]^and_result107[195]^and_result107[196]^and_result107[197]^and_result107[198]^and_result107[199]^and_result107[200]^and_result107[201]^and_result107[202]^and_result107[203]^and_result107[204]^and_result107[205]^and_result107[206]^and_result107[207]^and_result107[208]^and_result107[209]^and_result107[210]^and_result107[211]^and_result107[212]^and_result107[213]^and_result107[214]^and_result107[215]^and_result107[216]^and_result107[217]^and_result107[218]^and_result107[219]^and_result107[220]^and_result107[221]^and_result107[222]^and_result107[223]^and_result107[224]^and_result107[225]^and_result107[226]^and_result107[227]^and_result107[228]^and_result107[229]^and_result107[230]^and_result107[231]^and_result107[232]^and_result107[233]^and_result107[234]^and_result107[235]^and_result107[236]^and_result107[237]^and_result107[238]^and_result107[239]^and_result107[240]^and_result107[241]^and_result107[242]^and_result107[243]^and_result107[244]^and_result107[245]^and_result107[246]^and_result107[247]^and_result107[248]^and_result107[249]^and_result107[250]^and_result107[251]^and_result107[252]^and_result107[253]^and_result107[254];
assign key[108]=and_result108[0]^and_result108[1]^and_result108[2]^and_result108[3]^and_result108[4]^and_result108[5]^and_result108[6]^and_result108[7]^and_result108[8]^and_result108[9]^and_result108[10]^and_result108[11]^and_result108[12]^and_result108[13]^and_result108[14]^and_result108[15]^and_result108[16]^and_result108[17]^and_result108[18]^and_result108[19]^and_result108[20]^and_result108[21]^and_result108[22]^and_result108[23]^and_result108[24]^and_result108[25]^and_result108[26]^and_result108[27]^and_result108[28]^and_result108[29]^and_result108[30]^and_result108[31]^and_result108[32]^and_result108[33]^and_result108[34]^and_result108[35]^and_result108[36]^and_result108[37]^and_result108[38]^and_result108[39]^and_result108[40]^and_result108[41]^and_result108[42]^and_result108[43]^and_result108[44]^and_result108[45]^and_result108[46]^and_result108[47]^and_result108[48]^and_result108[49]^and_result108[50]^and_result108[51]^and_result108[52]^and_result108[53]^and_result108[54]^and_result108[55]^and_result108[56]^and_result108[57]^and_result108[58]^and_result108[59]^and_result108[60]^and_result108[61]^and_result108[62]^and_result108[63]^and_result108[64]^and_result108[65]^and_result108[66]^and_result108[67]^and_result108[68]^and_result108[69]^and_result108[70]^and_result108[71]^and_result108[72]^and_result108[73]^and_result108[74]^and_result108[75]^and_result108[76]^and_result108[77]^and_result108[78]^and_result108[79]^and_result108[80]^and_result108[81]^and_result108[82]^and_result108[83]^and_result108[84]^and_result108[85]^and_result108[86]^and_result108[87]^and_result108[88]^and_result108[89]^and_result108[90]^and_result108[91]^and_result108[92]^and_result108[93]^and_result108[94]^and_result108[95]^and_result108[96]^and_result108[97]^and_result108[98]^and_result108[99]^and_result108[100]^and_result108[101]^and_result108[102]^and_result108[103]^and_result108[104]^and_result108[105]^and_result108[106]^and_result108[107]^and_result108[108]^and_result108[109]^and_result108[110]^and_result108[111]^and_result108[112]^and_result108[113]^and_result108[114]^and_result108[115]^and_result108[116]^and_result108[117]^and_result108[118]^and_result108[119]^and_result108[120]^and_result108[121]^and_result108[122]^and_result108[123]^and_result108[124]^and_result108[125]^and_result108[126]^and_result108[127]^and_result108[128]^and_result108[129]^and_result108[130]^and_result108[131]^and_result108[132]^and_result108[133]^and_result108[134]^and_result108[135]^and_result108[136]^and_result108[137]^and_result108[138]^and_result108[139]^and_result108[140]^and_result108[141]^and_result108[142]^and_result108[143]^and_result108[144]^and_result108[145]^and_result108[146]^and_result108[147]^and_result108[148]^and_result108[149]^and_result108[150]^and_result108[151]^and_result108[152]^and_result108[153]^and_result108[154]^and_result108[155]^and_result108[156]^and_result108[157]^and_result108[158]^and_result108[159]^and_result108[160]^and_result108[161]^and_result108[162]^and_result108[163]^and_result108[164]^and_result108[165]^and_result108[166]^and_result108[167]^and_result108[168]^and_result108[169]^and_result108[170]^and_result108[171]^and_result108[172]^and_result108[173]^and_result108[174]^and_result108[175]^and_result108[176]^and_result108[177]^and_result108[178]^and_result108[179]^and_result108[180]^and_result108[181]^and_result108[182]^and_result108[183]^and_result108[184]^and_result108[185]^and_result108[186]^and_result108[187]^and_result108[188]^and_result108[189]^and_result108[190]^and_result108[191]^and_result108[192]^and_result108[193]^and_result108[194]^and_result108[195]^and_result108[196]^and_result108[197]^and_result108[198]^and_result108[199]^and_result108[200]^and_result108[201]^and_result108[202]^and_result108[203]^and_result108[204]^and_result108[205]^and_result108[206]^and_result108[207]^and_result108[208]^and_result108[209]^and_result108[210]^and_result108[211]^and_result108[212]^and_result108[213]^and_result108[214]^and_result108[215]^and_result108[216]^and_result108[217]^and_result108[218]^and_result108[219]^and_result108[220]^and_result108[221]^and_result108[222]^and_result108[223]^and_result108[224]^and_result108[225]^and_result108[226]^and_result108[227]^and_result108[228]^and_result108[229]^and_result108[230]^and_result108[231]^and_result108[232]^and_result108[233]^and_result108[234]^and_result108[235]^and_result108[236]^and_result108[237]^and_result108[238]^and_result108[239]^and_result108[240]^and_result108[241]^and_result108[242]^and_result108[243]^and_result108[244]^and_result108[245]^and_result108[246]^and_result108[247]^and_result108[248]^and_result108[249]^and_result108[250]^and_result108[251]^and_result108[252]^and_result108[253]^and_result108[254];
assign key[109]=and_result109[0]^and_result109[1]^and_result109[2]^and_result109[3]^and_result109[4]^and_result109[5]^and_result109[6]^and_result109[7]^and_result109[8]^and_result109[9]^and_result109[10]^and_result109[11]^and_result109[12]^and_result109[13]^and_result109[14]^and_result109[15]^and_result109[16]^and_result109[17]^and_result109[18]^and_result109[19]^and_result109[20]^and_result109[21]^and_result109[22]^and_result109[23]^and_result109[24]^and_result109[25]^and_result109[26]^and_result109[27]^and_result109[28]^and_result109[29]^and_result109[30]^and_result109[31]^and_result109[32]^and_result109[33]^and_result109[34]^and_result109[35]^and_result109[36]^and_result109[37]^and_result109[38]^and_result109[39]^and_result109[40]^and_result109[41]^and_result109[42]^and_result109[43]^and_result109[44]^and_result109[45]^and_result109[46]^and_result109[47]^and_result109[48]^and_result109[49]^and_result109[50]^and_result109[51]^and_result109[52]^and_result109[53]^and_result109[54]^and_result109[55]^and_result109[56]^and_result109[57]^and_result109[58]^and_result109[59]^and_result109[60]^and_result109[61]^and_result109[62]^and_result109[63]^and_result109[64]^and_result109[65]^and_result109[66]^and_result109[67]^and_result109[68]^and_result109[69]^and_result109[70]^and_result109[71]^and_result109[72]^and_result109[73]^and_result109[74]^and_result109[75]^and_result109[76]^and_result109[77]^and_result109[78]^and_result109[79]^and_result109[80]^and_result109[81]^and_result109[82]^and_result109[83]^and_result109[84]^and_result109[85]^and_result109[86]^and_result109[87]^and_result109[88]^and_result109[89]^and_result109[90]^and_result109[91]^and_result109[92]^and_result109[93]^and_result109[94]^and_result109[95]^and_result109[96]^and_result109[97]^and_result109[98]^and_result109[99]^and_result109[100]^and_result109[101]^and_result109[102]^and_result109[103]^and_result109[104]^and_result109[105]^and_result109[106]^and_result109[107]^and_result109[108]^and_result109[109]^and_result109[110]^and_result109[111]^and_result109[112]^and_result109[113]^and_result109[114]^and_result109[115]^and_result109[116]^and_result109[117]^and_result109[118]^and_result109[119]^and_result109[120]^and_result109[121]^and_result109[122]^and_result109[123]^and_result109[124]^and_result109[125]^and_result109[126]^and_result109[127]^and_result109[128]^and_result109[129]^and_result109[130]^and_result109[131]^and_result109[132]^and_result109[133]^and_result109[134]^and_result109[135]^and_result109[136]^and_result109[137]^and_result109[138]^and_result109[139]^and_result109[140]^and_result109[141]^and_result109[142]^and_result109[143]^and_result109[144]^and_result109[145]^and_result109[146]^and_result109[147]^and_result109[148]^and_result109[149]^and_result109[150]^and_result109[151]^and_result109[152]^and_result109[153]^and_result109[154]^and_result109[155]^and_result109[156]^and_result109[157]^and_result109[158]^and_result109[159]^and_result109[160]^and_result109[161]^and_result109[162]^and_result109[163]^and_result109[164]^and_result109[165]^and_result109[166]^and_result109[167]^and_result109[168]^and_result109[169]^and_result109[170]^and_result109[171]^and_result109[172]^and_result109[173]^and_result109[174]^and_result109[175]^and_result109[176]^and_result109[177]^and_result109[178]^and_result109[179]^and_result109[180]^and_result109[181]^and_result109[182]^and_result109[183]^and_result109[184]^and_result109[185]^and_result109[186]^and_result109[187]^and_result109[188]^and_result109[189]^and_result109[190]^and_result109[191]^and_result109[192]^and_result109[193]^and_result109[194]^and_result109[195]^and_result109[196]^and_result109[197]^and_result109[198]^and_result109[199]^and_result109[200]^and_result109[201]^and_result109[202]^and_result109[203]^and_result109[204]^and_result109[205]^and_result109[206]^and_result109[207]^and_result109[208]^and_result109[209]^and_result109[210]^and_result109[211]^and_result109[212]^and_result109[213]^and_result109[214]^and_result109[215]^and_result109[216]^and_result109[217]^and_result109[218]^and_result109[219]^and_result109[220]^and_result109[221]^and_result109[222]^and_result109[223]^and_result109[224]^and_result109[225]^and_result109[226]^and_result109[227]^and_result109[228]^and_result109[229]^and_result109[230]^and_result109[231]^and_result109[232]^and_result109[233]^and_result109[234]^and_result109[235]^and_result109[236]^and_result109[237]^and_result109[238]^and_result109[239]^and_result109[240]^and_result109[241]^and_result109[242]^and_result109[243]^and_result109[244]^and_result109[245]^and_result109[246]^and_result109[247]^and_result109[248]^and_result109[249]^and_result109[250]^and_result109[251]^and_result109[252]^and_result109[253]^and_result109[254];
assign key[110]=and_result110[0]^and_result110[1]^and_result110[2]^and_result110[3]^and_result110[4]^and_result110[5]^and_result110[6]^and_result110[7]^and_result110[8]^and_result110[9]^and_result110[10]^and_result110[11]^and_result110[12]^and_result110[13]^and_result110[14]^and_result110[15]^and_result110[16]^and_result110[17]^and_result110[18]^and_result110[19]^and_result110[20]^and_result110[21]^and_result110[22]^and_result110[23]^and_result110[24]^and_result110[25]^and_result110[26]^and_result110[27]^and_result110[28]^and_result110[29]^and_result110[30]^and_result110[31]^and_result110[32]^and_result110[33]^and_result110[34]^and_result110[35]^and_result110[36]^and_result110[37]^and_result110[38]^and_result110[39]^and_result110[40]^and_result110[41]^and_result110[42]^and_result110[43]^and_result110[44]^and_result110[45]^and_result110[46]^and_result110[47]^and_result110[48]^and_result110[49]^and_result110[50]^and_result110[51]^and_result110[52]^and_result110[53]^and_result110[54]^and_result110[55]^and_result110[56]^and_result110[57]^and_result110[58]^and_result110[59]^and_result110[60]^and_result110[61]^and_result110[62]^and_result110[63]^and_result110[64]^and_result110[65]^and_result110[66]^and_result110[67]^and_result110[68]^and_result110[69]^and_result110[70]^and_result110[71]^and_result110[72]^and_result110[73]^and_result110[74]^and_result110[75]^and_result110[76]^and_result110[77]^and_result110[78]^and_result110[79]^and_result110[80]^and_result110[81]^and_result110[82]^and_result110[83]^and_result110[84]^and_result110[85]^and_result110[86]^and_result110[87]^and_result110[88]^and_result110[89]^and_result110[90]^and_result110[91]^and_result110[92]^and_result110[93]^and_result110[94]^and_result110[95]^and_result110[96]^and_result110[97]^and_result110[98]^and_result110[99]^and_result110[100]^and_result110[101]^and_result110[102]^and_result110[103]^and_result110[104]^and_result110[105]^and_result110[106]^and_result110[107]^and_result110[108]^and_result110[109]^and_result110[110]^and_result110[111]^and_result110[112]^and_result110[113]^and_result110[114]^and_result110[115]^and_result110[116]^and_result110[117]^and_result110[118]^and_result110[119]^and_result110[120]^and_result110[121]^and_result110[122]^and_result110[123]^and_result110[124]^and_result110[125]^and_result110[126]^and_result110[127]^and_result110[128]^and_result110[129]^and_result110[130]^and_result110[131]^and_result110[132]^and_result110[133]^and_result110[134]^and_result110[135]^and_result110[136]^and_result110[137]^and_result110[138]^and_result110[139]^and_result110[140]^and_result110[141]^and_result110[142]^and_result110[143]^and_result110[144]^and_result110[145]^and_result110[146]^and_result110[147]^and_result110[148]^and_result110[149]^and_result110[150]^and_result110[151]^and_result110[152]^and_result110[153]^and_result110[154]^and_result110[155]^and_result110[156]^and_result110[157]^and_result110[158]^and_result110[159]^and_result110[160]^and_result110[161]^and_result110[162]^and_result110[163]^and_result110[164]^and_result110[165]^and_result110[166]^and_result110[167]^and_result110[168]^and_result110[169]^and_result110[170]^and_result110[171]^and_result110[172]^and_result110[173]^and_result110[174]^and_result110[175]^and_result110[176]^and_result110[177]^and_result110[178]^and_result110[179]^and_result110[180]^and_result110[181]^and_result110[182]^and_result110[183]^and_result110[184]^and_result110[185]^and_result110[186]^and_result110[187]^and_result110[188]^and_result110[189]^and_result110[190]^and_result110[191]^and_result110[192]^and_result110[193]^and_result110[194]^and_result110[195]^and_result110[196]^and_result110[197]^and_result110[198]^and_result110[199]^and_result110[200]^and_result110[201]^and_result110[202]^and_result110[203]^and_result110[204]^and_result110[205]^and_result110[206]^and_result110[207]^and_result110[208]^and_result110[209]^and_result110[210]^and_result110[211]^and_result110[212]^and_result110[213]^and_result110[214]^and_result110[215]^and_result110[216]^and_result110[217]^and_result110[218]^and_result110[219]^and_result110[220]^and_result110[221]^and_result110[222]^and_result110[223]^and_result110[224]^and_result110[225]^and_result110[226]^and_result110[227]^and_result110[228]^and_result110[229]^and_result110[230]^and_result110[231]^and_result110[232]^and_result110[233]^and_result110[234]^and_result110[235]^and_result110[236]^and_result110[237]^and_result110[238]^and_result110[239]^and_result110[240]^and_result110[241]^and_result110[242]^and_result110[243]^and_result110[244]^and_result110[245]^and_result110[246]^and_result110[247]^and_result110[248]^and_result110[249]^and_result110[250]^and_result110[251]^and_result110[252]^and_result110[253]^and_result110[254];
assign key[111]=and_result111[0]^and_result111[1]^and_result111[2]^and_result111[3]^and_result111[4]^and_result111[5]^and_result111[6]^and_result111[7]^and_result111[8]^and_result111[9]^and_result111[10]^and_result111[11]^and_result111[12]^and_result111[13]^and_result111[14]^and_result111[15]^and_result111[16]^and_result111[17]^and_result111[18]^and_result111[19]^and_result111[20]^and_result111[21]^and_result111[22]^and_result111[23]^and_result111[24]^and_result111[25]^and_result111[26]^and_result111[27]^and_result111[28]^and_result111[29]^and_result111[30]^and_result111[31]^and_result111[32]^and_result111[33]^and_result111[34]^and_result111[35]^and_result111[36]^and_result111[37]^and_result111[38]^and_result111[39]^and_result111[40]^and_result111[41]^and_result111[42]^and_result111[43]^and_result111[44]^and_result111[45]^and_result111[46]^and_result111[47]^and_result111[48]^and_result111[49]^and_result111[50]^and_result111[51]^and_result111[52]^and_result111[53]^and_result111[54]^and_result111[55]^and_result111[56]^and_result111[57]^and_result111[58]^and_result111[59]^and_result111[60]^and_result111[61]^and_result111[62]^and_result111[63]^and_result111[64]^and_result111[65]^and_result111[66]^and_result111[67]^and_result111[68]^and_result111[69]^and_result111[70]^and_result111[71]^and_result111[72]^and_result111[73]^and_result111[74]^and_result111[75]^and_result111[76]^and_result111[77]^and_result111[78]^and_result111[79]^and_result111[80]^and_result111[81]^and_result111[82]^and_result111[83]^and_result111[84]^and_result111[85]^and_result111[86]^and_result111[87]^and_result111[88]^and_result111[89]^and_result111[90]^and_result111[91]^and_result111[92]^and_result111[93]^and_result111[94]^and_result111[95]^and_result111[96]^and_result111[97]^and_result111[98]^and_result111[99]^and_result111[100]^and_result111[101]^and_result111[102]^and_result111[103]^and_result111[104]^and_result111[105]^and_result111[106]^and_result111[107]^and_result111[108]^and_result111[109]^and_result111[110]^and_result111[111]^and_result111[112]^and_result111[113]^and_result111[114]^and_result111[115]^and_result111[116]^and_result111[117]^and_result111[118]^and_result111[119]^and_result111[120]^and_result111[121]^and_result111[122]^and_result111[123]^and_result111[124]^and_result111[125]^and_result111[126]^and_result111[127]^and_result111[128]^and_result111[129]^and_result111[130]^and_result111[131]^and_result111[132]^and_result111[133]^and_result111[134]^and_result111[135]^and_result111[136]^and_result111[137]^and_result111[138]^and_result111[139]^and_result111[140]^and_result111[141]^and_result111[142]^and_result111[143]^and_result111[144]^and_result111[145]^and_result111[146]^and_result111[147]^and_result111[148]^and_result111[149]^and_result111[150]^and_result111[151]^and_result111[152]^and_result111[153]^and_result111[154]^and_result111[155]^and_result111[156]^and_result111[157]^and_result111[158]^and_result111[159]^and_result111[160]^and_result111[161]^and_result111[162]^and_result111[163]^and_result111[164]^and_result111[165]^and_result111[166]^and_result111[167]^and_result111[168]^and_result111[169]^and_result111[170]^and_result111[171]^and_result111[172]^and_result111[173]^and_result111[174]^and_result111[175]^and_result111[176]^and_result111[177]^and_result111[178]^and_result111[179]^and_result111[180]^and_result111[181]^and_result111[182]^and_result111[183]^and_result111[184]^and_result111[185]^and_result111[186]^and_result111[187]^and_result111[188]^and_result111[189]^and_result111[190]^and_result111[191]^and_result111[192]^and_result111[193]^and_result111[194]^and_result111[195]^and_result111[196]^and_result111[197]^and_result111[198]^and_result111[199]^and_result111[200]^and_result111[201]^and_result111[202]^and_result111[203]^and_result111[204]^and_result111[205]^and_result111[206]^and_result111[207]^and_result111[208]^and_result111[209]^and_result111[210]^and_result111[211]^and_result111[212]^and_result111[213]^and_result111[214]^and_result111[215]^and_result111[216]^and_result111[217]^and_result111[218]^and_result111[219]^and_result111[220]^and_result111[221]^and_result111[222]^and_result111[223]^and_result111[224]^and_result111[225]^and_result111[226]^and_result111[227]^and_result111[228]^and_result111[229]^and_result111[230]^and_result111[231]^and_result111[232]^and_result111[233]^and_result111[234]^and_result111[235]^and_result111[236]^and_result111[237]^and_result111[238]^and_result111[239]^and_result111[240]^and_result111[241]^and_result111[242]^and_result111[243]^and_result111[244]^and_result111[245]^and_result111[246]^and_result111[247]^and_result111[248]^and_result111[249]^and_result111[250]^and_result111[251]^and_result111[252]^and_result111[253]^and_result111[254];
assign key[112]=and_result112[0]^and_result112[1]^and_result112[2]^and_result112[3]^and_result112[4]^and_result112[5]^and_result112[6]^and_result112[7]^and_result112[8]^and_result112[9]^and_result112[10]^and_result112[11]^and_result112[12]^and_result112[13]^and_result112[14]^and_result112[15]^and_result112[16]^and_result112[17]^and_result112[18]^and_result112[19]^and_result112[20]^and_result112[21]^and_result112[22]^and_result112[23]^and_result112[24]^and_result112[25]^and_result112[26]^and_result112[27]^and_result112[28]^and_result112[29]^and_result112[30]^and_result112[31]^and_result112[32]^and_result112[33]^and_result112[34]^and_result112[35]^and_result112[36]^and_result112[37]^and_result112[38]^and_result112[39]^and_result112[40]^and_result112[41]^and_result112[42]^and_result112[43]^and_result112[44]^and_result112[45]^and_result112[46]^and_result112[47]^and_result112[48]^and_result112[49]^and_result112[50]^and_result112[51]^and_result112[52]^and_result112[53]^and_result112[54]^and_result112[55]^and_result112[56]^and_result112[57]^and_result112[58]^and_result112[59]^and_result112[60]^and_result112[61]^and_result112[62]^and_result112[63]^and_result112[64]^and_result112[65]^and_result112[66]^and_result112[67]^and_result112[68]^and_result112[69]^and_result112[70]^and_result112[71]^and_result112[72]^and_result112[73]^and_result112[74]^and_result112[75]^and_result112[76]^and_result112[77]^and_result112[78]^and_result112[79]^and_result112[80]^and_result112[81]^and_result112[82]^and_result112[83]^and_result112[84]^and_result112[85]^and_result112[86]^and_result112[87]^and_result112[88]^and_result112[89]^and_result112[90]^and_result112[91]^and_result112[92]^and_result112[93]^and_result112[94]^and_result112[95]^and_result112[96]^and_result112[97]^and_result112[98]^and_result112[99]^and_result112[100]^and_result112[101]^and_result112[102]^and_result112[103]^and_result112[104]^and_result112[105]^and_result112[106]^and_result112[107]^and_result112[108]^and_result112[109]^and_result112[110]^and_result112[111]^and_result112[112]^and_result112[113]^and_result112[114]^and_result112[115]^and_result112[116]^and_result112[117]^and_result112[118]^and_result112[119]^and_result112[120]^and_result112[121]^and_result112[122]^and_result112[123]^and_result112[124]^and_result112[125]^and_result112[126]^and_result112[127]^and_result112[128]^and_result112[129]^and_result112[130]^and_result112[131]^and_result112[132]^and_result112[133]^and_result112[134]^and_result112[135]^and_result112[136]^and_result112[137]^and_result112[138]^and_result112[139]^and_result112[140]^and_result112[141]^and_result112[142]^and_result112[143]^and_result112[144]^and_result112[145]^and_result112[146]^and_result112[147]^and_result112[148]^and_result112[149]^and_result112[150]^and_result112[151]^and_result112[152]^and_result112[153]^and_result112[154]^and_result112[155]^and_result112[156]^and_result112[157]^and_result112[158]^and_result112[159]^and_result112[160]^and_result112[161]^and_result112[162]^and_result112[163]^and_result112[164]^and_result112[165]^and_result112[166]^and_result112[167]^and_result112[168]^and_result112[169]^and_result112[170]^and_result112[171]^and_result112[172]^and_result112[173]^and_result112[174]^and_result112[175]^and_result112[176]^and_result112[177]^and_result112[178]^and_result112[179]^and_result112[180]^and_result112[181]^and_result112[182]^and_result112[183]^and_result112[184]^and_result112[185]^and_result112[186]^and_result112[187]^and_result112[188]^and_result112[189]^and_result112[190]^and_result112[191]^and_result112[192]^and_result112[193]^and_result112[194]^and_result112[195]^and_result112[196]^and_result112[197]^and_result112[198]^and_result112[199]^and_result112[200]^and_result112[201]^and_result112[202]^and_result112[203]^and_result112[204]^and_result112[205]^and_result112[206]^and_result112[207]^and_result112[208]^and_result112[209]^and_result112[210]^and_result112[211]^and_result112[212]^and_result112[213]^and_result112[214]^and_result112[215]^and_result112[216]^and_result112[217]^and_result112[218]^and_result112[219]^and_result112[220]^and_result112[221]^and_result112[222]^and_result112[223]^and_result112[224]^and_result112[225]^and_result112[226]^and_result112[227]^and_result112[228]^and_result112[229]^and_result112[230]^and_result112[231]^and_result112[232]^and_result112[233]^and_result112[234]^and_result112[235]^and_result112[236]^and_result112[237]^and_result112[238]^and_result112[239]^and_result112[240]^and_result112[241]^and_result112[242]^and_result112[243]^and_result112[244]^and_result112[245]^and_result112[246]^and_result112[247]^and_result112[248]^and_result112[249]^and_result112[250]^and_result112[251]^and_result112[252]^and_result112[253]^and_result112[254];
assign key[113]=and_result113[0]^and_result113[1]^and_result113[2]^and_result113[3]^and_result113[4]^and_result113[5]^and_result113[6]^and_result113[7]^and_result113[8]^and_result113[9]^and_result113[10]^and_result113[11]^and_result113[12]^and_result113[13]^and_result113[14]^and_result113[15]^and_result113[16]^and_result113[17]^and_result113[18]^and_result113[19]^and_result113[20]^and_result113[21]^and_result113[22]^and_result113[23]^and_result113[24]^and_result113[25]^and_result113[26]^and_result113[27]^and_result113[28]^and_result113[29]^and_result113[30]^and_result113[31]^and_result113[32]^and_result113[33]^and_result113[34]^and_result113[35]^and_result113[36]^and_result113[37]^and_result113[38]^and_result113[39]^and_result113[40]^and_result113[41]^and_result113[42]^and_result113[43]^and_result113[44]^and_result113[45]^and_result113[46]^and_result113[47]^and_result113[48]^and_result113[49]^and_result113[50]^and_result113[51]^and_result113[52]^and_result113[53]^and_result113[54]^and_result113[55]^and_result113[56]^and_result113[57]^and_result113[58]^and_result113[59]^and_result113[60]^and_result113[61]^and_result113[62]^and_result113[63]^and_result113[64]^and_result113[65]^and_result113[66]^and_result113[67]^and_result113[68]^and_result113[69]^and_result113[70]^and_result113[71]^and_result113[72]^and_result113[73]^and_result113[74]^and_result113[75]^and_result113[76]^and_result113[77]^and_result113[78]^and_result113[79]^and_result113[80]^and_result113[81]^and_result113[82]^and_result113[83]^and_result113[84]^and_result113[85]^and_result113[86]^and_result113[87]^and_result113[88]^and_result113[89]^and_result113[90]^and_result113[91]^and_result113[92]^and_result113[93]^and_result113[94]^and_result113[95]^and_result113[96]^and_result113[97]^and_result113[98]^and_result113[99]^and_result113[100]^and_result113[101]^and_result113[102]^and_result113[103]^and_result113[104]^and_result113[105]^and_result113[106]^and_result113[107]^and_result113[108]^and_result113[109]^and_result113[110]^and_result113[111]^and_result113[112]^and_result113[113]^and_result113[114]^and_result113[115]^and_result113[116]^and_result113[117]^and_result113[118]^and_result113[119]^and_result113[120]^and_result113[121]^and_result113[122]^and_result113[123]^and_result113[124]^and_result113[125]^and_result113[126]^and_result113[127]^and_result113[128]^and_result113[129]^and_result113[130]^and_result113[131]^and_result113[132]^and_result113[133]^and_result113[134]^and_result113[135]^and_result113[136]^and_result113[137]^and_result113[138]^and_result113[139]^and_result113[140]^and_result113[141]^and_result113[142]^and_result113[143]^and_result113[144]^and_result113[145]^and_result113[146]^and_result113[147]^and_result113[148]^and_result113[149]^and_result113[150]^and_result113[151]^and_result113[152]^and_result113[153]^and_result113[154]^and_result113[155]^and_result113[156]^and_result113[157]^and_result113[158]^and_result113[159]^and_result113[160]^and_result113[161]^and_result113[162]^and_result113[163]^and_result113[164]^and_result113[165]^and_result113[166]^and_result113[167]^and_result113[168]^and_result113[169]^and_result113[170]^and_result113[171]^and_result113[172]^and_result113[173]^and_result113[174]^and_result113[175]^and_result113[176]^and_result113[177]^and_result113[178]^and_result113[179]^and_result113[180]^and_result113[181]^and_result113[182]^and_result113[183]^and_result113[184]^and_result113[185]^and_result113[186]^and_result113[187]^and_result113[188]^and_result113[189]^and_result113[190]^and_result113[191]^and_result113[192]^and_result113[193]^and_result113[194]^and_result113[195]^and_result113[196]^and_result113[197]^and_result113[198]^and_result113[199]^and_result113[200]^and_result113[201]^and_result113[202]^and_result113[203]^and_result113[204]^and_result113[205]^and_result113[206]^and_result113[207]^and_result113[208]^and_result113[209]^and_result113[210]^and_result113[211]^and_result113[212]^and_result113[213]^and_result113[214]^and_result113[215]^and_result113[216]^and_result113[217]^and_result113[218]^and_result113[219]^and_result113[220]^and_result113[221]^and_result113[222]^and_result113[223]^and_result113[224]^and_result113[225]^and_result113[226]^and_result113[227]^and_result113[228]^and_result113[229]^and_result113[230]^and_result113[231]^and_result113[232]^and_result113[233]^and_result113[234]^and_result113[235]^and_result113[236]^and_result113[237]^and_result113[238]^and_result113[239]^and_result113[240]^and_result113[241]^and_result113[242]^and_result113[243]^and_result113[244]^and_result113[245]^and_result113[246]^and_result113[247]^and_result113[248]^and_result113[249]^and_result113[250]^and_result113[251]^and_result113[252]^and_result113[253]^and_result113[254];
assign key[114]=and_result114[0]^and_result114[1]^and_result114[2]^and_result114[3]^and_result114[4]^and_result114[5]^and_result114[6]^and_result114[7]^and_result114[8]^and_result114[9]^and_result114[10]^and_result114[11]^and_result114[12]^and_result114[13]^and_result114[14]^and_result114[15]^and_result114[16]^and_result114[17]^and_result114[18]^and_result114[19]^and_result114[20]^and_result114[21]^and_result114[22]^and_result114[23]^and_result114[24]^and_result114[25]^and_result114[26]^and_result114[27]^and_result114[28]^and_result114[29]^and_result114[30]^and_result114[31]^and_result114[32]^and_result114[33]^and_result114[34]^and_result114[35]^and_result114[36]^and_result114[37]^and_result114[38]^and_result114[39]^and_result114[40]^and_result114[41]^and_result114[42]^and_result114[43]^and_result114[44]^and_result114[45]^and_result114[46]^and_result114[47]^and_result114[48]^and_result114[49]^and_result114[50]^and_result114[51]^and_result114[52]^and_result114[53]^and_result114[54]^and_result114[55]^and_result114[56]^and_result114[57]^and_result114[58]^and_result114[59]^and_result114[60]^and_result114[61]^and_result114[62]^and_result114[63]^and_result114[64]^and_result114[65]^and_result114[66]^and_result114[67]^and_result114[68]^and_result114[69]^and_result114[70]^and_result114[71]^and_result114[72]^and_result114[73]^and_result114[74]^and_result114[75]^and_result114[76]^and_result114[77]^and_result114[78]^and_result114[79]^and_result114[80]^and_result114[81]^and_result114[82]^and_result114[83]^and_result114[84]^and_result114[85]^and_result114[86]^and_result114[87]^and_result114[88]^and_result114[89]^and_result114[90]^and_result114[91]^and_result114[92]^and_result114[93]^and_result114[94]^and_result114[95]^and_result114[96]^and_result114[97]^and_result114[98]^and_result114[99]^and_result114[100]^and_result114[101]^and_result114[102]^and_result114[103]^and_result114[104]^and_result114[105]^and_result114[106]^and_result114[107]^and_result114[108]^and_result114[109]^and_result114[110]^and_result114[111]^and_result114[112]^and_result114[113]^and_result114[114]^and_result114[115]^and_result114[116]^and_result114[117]^and_result114[118]^and_result114[119]^and_result114[120]^and_result114[121]^and_result114[122]^and_result114[123]^and_result114[124]^and_result114[125]^and_result114[126]^and_result114[127]^and_result114[128]^and_result114[129]^and_result114[130]^and_result114[131]^and_result114[132]^and_result114[133]^and_result114[134]^and_result114[135]^and_result114[136]^and_result114[137]^and_result114[138]^and_result114[139]^and_result114[140]^and_result114[141]^and_result114[142]^and_result114[143]^and_result114[144]^and_result114[145]^and_result114[146]^and_result114[147]^and_result114[148]^and_result114[149]^and_result114[150]^and_result114[151]^and_result114[152]^and_result114[153]^and_result114[154]^and_result114[155]^and_result114[156]^and_result114[157]^and_result114[158]^and_result114[159]^and_result114[160]^and_result114[161]^and_result114[162]^and_result114[163]^and_result114[164]^and_result114[165]^and_result114[166]^and_result114[167]^and_result114[168]^and_result114[169]^and_result114[170]^and_result114[171]^and_result114[172]^and_result114[173]^and_result114[174]^and_result114[175]^and_result114[176]^and_result114[177]^and_result114[178]^and_result114[179]^and_result114[180]^and_result114[181]^and_result114[182]^and_result114[183]^and_result114[184]^and_result114[185]^and_result114[186]^and_result114[187]^and_result114[188]^and_result114[189]^and_result114[190]^and_result114[191]^and_result114[192]^and_result114[193]^and_result114[194]^and_result114[195]^and_result114[196]^and_result114[197]^and_result114[198]^and_result114[199]^and_result114[200]^and_result114[201]^and_result114[202]^and_result114[203]^and_result114[204]^and_result114[205]^and_result114[206]^and_result114[207]^and_result114[208]^and_result114[209]^and_result114[210]^and_result114[211]^and_result114[212]^and_result114[213]^and_result114[214]^and_result114[215]^and_result114[216]^and_result114[217]^and_result114[218]^and_result114[219]^and_result114[220]^and_result114[221]^and_result114[222]^and_result114[223]^and_result114[224]^and_result114[225]^and_result114[226]^and_result114[227]^and_result114[228]^and_result114[229]^and_result114[230]^and_result114[231]^and_result114[232]^and_result114[233]^and_result114[234]^and_result114[235]^and_result114[236]^and_result114[237]^and_result114[238]^and_result114[239]^and_result114[240]^and_result114[241]^and_result114[242]^and_result114[243]^and_result114[244]^and_result114[245]^and_result114[246]^and_result114[247]^and_result114[248]^and_result114[249]^and_result114[250]^and_result114[251]^and_result114[252]^and_result114[253]^and_result114[254];
assign key[115]=and_result115[0]^and_result115[1]^and_result115[2]^and_result115[3]^and_result115[4]^and_result115[5]^and_result115[6]^and_result115[7]^and_result115[8]^and_result115[9]^and_result115[10]^and_result115[11]^and_result115[12]^and_result115[13]^and_result115[14]^and_result115[15]^and_result115[16]^and_result115[17]^and_result115[18]^and_result115[19]^and_result115[20]^and_result115[21]^and_result115[22]^and_result115[23]^and_result115[24]^and_result115[25]^and_result115[26]^and_result115[27]^and_result115[28]^and_result115[29]^and_result115[30]^and_result115[31]^and_result115[32]^and_result115[33]^and_result115[34]^and_result115[35]^and_result115[36]^and_result115[37]^and_result115[38]^and_result115[39]^and_result115[40]^and_result115[41]^and_result115[42]^and_result115[43]^and_result115[44]^and_result115[45]^and_result115[46]^and_result115[47]^and_result115[48]^and_result115[49]^and_result115[50]^and_result115[51]^and_result115[52]^and_result115[53]^and_result115[54]^and_result115[55]^and_result115[56]^and_result115[57]^and_result115[58]^and_result115[59]^and_result115[60]^and_result115[61]^and_result115[62]^and_result115[63]^and_result115[64]^and_result115[65]^and_result115[66]^and_result115[67]^and_result115[68]^and_result115[69]^and_result115[70]^and_result115[71]^and_result115[72]^and_result115[73]^and_result115[74]^and_result115[75]^and_result115[76]^and_result115[77]^and_result115[78]^and_result115[79]^and_result115[80]^and_result115[81]^and_result115[82]^and_result115[83]^and_result115[84]^and_result115[85]^and_result115[86]^and_result115[87]^and_result115[88]^and_result115[89]^and_result115[90]^and_result115[91]^and_result115[92]^and_result115[93]^and_result115[94]^and_result115[95]^and_result115[96]^and_result115[97]^and_result115[98]^and_result115[99]^and_result115[100]^and_result115[101]^and_result115[102]^and_result115[103]^and_result115[104]^and_result115[105]^and_result115[106]^and_result115[107]^and_result115[108]^and_result115[109]^and_result115[110]^and_result115[111]^and_result115[112]^and_result115[113]^and_result115[114]^and_result115[115]^and_result115[116]^and_result115[117]^and_result115[118]^and_result115[119]^and_result115[120]^and_result115[121]^and_result115[122]^and_result115[123]^and_result115[124]^and_result115[125]^and_result115[126]^and_result115[127]^and_result115[128]^and_result115[129]^and_result115[130]^and_result115[131]^and_result115[132]^and_result115[133]^and_result115[134]^and_result115[135]^and_result115[136]^and_result115[137]^and_result115[138]^and_result115[139]^and_result115[140]^and_result115[141]^and_result115[142]^and_result115[143]^and_result115[144]^and_result115[145]^and_result115[146]^and_result115[147]^and_result115[148]^and_result115[149]^and_result115[150]^and_result115[151]^and_result115[152]^and_result115[153]^and_result115[154]^and_result115[155]^and_result115[156]^and_result115[157]^and_result115[158]^and_result115[159]^and_result115[160]^and_result115[161]^and_result115[162]^and_result115[163]^and_result115[164]^and_result115[165]^and_result115[166]^and_result115[167]^and_result115[168]^and_result115[169]^and_result115[170]^and_result115[171]^and_result115[172]^and_result115[173]^and_result115[174]^and_result115[175]^and_result115[176]^and_result115[177]^and_result115[178]^and_result115[179]^and_result115[180]^and_result115[181]^and_result115[182]^and_result115[183]^and_result115[184]^and_result115[185]^and_result115[186]^and_result115[187]^and_result115[188]^and_result115[189]^and_result115[190]^and_result115[191]^and_result115[192]^and_result115[193]^and_result115[194]^and_result115[195]^and_result115[196]^and_result115[197]^and_result115[198]^and_result115[199]^and_result115[200]^and_result115[201]^and_result115[202]^and_result115[203]^and_result115[204]^and_result115[205]^and_result115[206]^and_result115[207]^and_result115[208]^and_result115[209]^and_result115[210]^and_result115[211]^and_result115[212]^and_result115[213]^and_result115[214]^and_result115[215]^and_result115[216]^and_result115[217]^and_result115[218]^and_result115[219]^and_result115[220]^and_result115[221]^and_result115[222]^and_result115[223]^and_result115[224]^and_result115[225]^and_result115[226]^and_result115[227]^and_result115[228]^and_result115[229]^and_result115[230]^and_result115[231]^and_result115[232]^and_result115[233]^and_result115[234]^and_result115[235]^and_result115[236]^and_result115[237]^and_result115[238]^and_result115[239]^and_result115[240]^and_result115[241]^and_result115[242]^and_result115[243]^and_result115[244]^and_result115[245]^and_result115[246]^and_result115[247]^and_result115[248]^and_result115[249]^and_result115[250]^and_result115[251]^and_result115[252]^and_result115[253]^and_result115[254];
assign key[116]=and_result116[0]^and_result116[1]^and_result116[2]^and_result116[3]^and_result116[4]^and_result116[5]^and_result116[6]^and_result116[7]^and_result116[8]^and_result116[9]^and_result116[10]^and_result116[11]^and_result116[12]^and_result116[13]^and_result116[14]^and_result116[15]^and_result116[16]^and_result116[17]^and_result116[18]^and_result116[19]^and_result116[20]^and_result116[21]^and_result116[22]^and_result116[23]^and_result116[24]^and_result116[25]^and_result116[26]^and_result116[27]^and_result116[28]^and_result116[29]^and_result116[30]^and_result116[31]^and_result116[32]^and_result116[33]^and_result116[34]^and_result116[35]^and_result116[36]^and_result116[37]^and_result116[38]^and_result116[39]^and_result116[40]^and_result116[41]^and_result116[42]^and_result116[43]^and_result116[44]^and_result116[45]^and_result116[46]^and_result116[47]^and_result116[48]^and_result116[49]^and_result116[50]^and_result116[51]^and_result116[52]^and_result116[53]^and_result116[54]^and_result116[55]^and_result116[56]^and_result116[57]^and_result116[58]^and_result116[59]^and_result116[60]^and_result116[61]^and_result116[62]^and_result116[63]^and_result116[64]^and_result116[65]^and_result116[66]^and_result116[67]^and_result116[68]^and_result116[69]^and_result116[70]^and_result116[71]^and_result116[72]^and_result116[73]^and_result116[74]^and_result116[75]^and_result116[76]^and_result116[77]^and_result116[78]^and_result116[79]^and_result116[80]^and_result116[81]^and_result116[82]^and_result116[83]^and_result116[84]^and_result116[85]^and_result116[86]^and_result116[87]^and_result116[88]^and_result116[89]^and_result116[90]^and_result116[91]^and_result116[92]^and_result116[93]^and_result116[94]^and_result116[95]^and_result116[96]^and_result116[97]^and_result116[98]^and_result116[99]^and_result116[100]^and_result116[101]^and_result116[102]^and_result116[103]^and_result116[104]^and_result116[105]^and_result116[106]^and_result116[107]^and_result116[108]^and_result116[109]^and_result116[110]^and_result116[111]^and_result116[112]^and_result116[113]^and_result116[114]^and_result116[115]^and_result116[116]^and_result116[117]^and_result116[118]^and_result116[119]^and_result116[120]^and_result116[121]^and_result116[122]^and_result116[123]^and_result116[124]^and_result116[125]^and_result116[126]^and_result116[127]^and_result116[128]^and_result116[129]^and_result116[130]^and_result116[131]^and_result116[132]^and_result116[133]^and_result116[134]^and_result116[135]^and_result116[136]^and_result116[137]^and_result116[138]^and_result116[139]^and_result116[140]^and_result116[141]^and_result116[142]^and_result116[143]^and_result116[144]^and_result116[145]^and_result116[146]^and_result116[147]^and_result116[148]^and_result116[149]^and_result116[150]^and_result116[151]^and_result116[152]^and_result116[153]^and_result116[154]^and_result116[155]^and_result116[156]^and_result116[157]^and_result116[158]^and_result116[159]^and_result116[160]^and_result116[161]^and_result116[162]^and_result116[163]^and_result116[164]^and_result116[165]^and_result116[166]^and_result116[167]^and_result116[168]^and_result116[169]^and_result116[170]^and_result116[171]^and_result116[172]^and_result116[173]^and_result116[174]^and_result116[175]^and_result116[176]^and_result116[177]^and_result116[178]^and_result116[179]^and_result116[180]^and_result116[181]^and_result116[182]^and_result116[183]^and_result116[184]^and_result116[185]^and_result116[186]^and_result116[187]^and_result116[188]^and_result116[189]^and_result116[190]^and_result116[191]^and_result116[192]^and_result116[193]^and_result116[194]^and_result116[195]^and_result116[196]^and_result116[197]^and_result116[198]^and_result116[199]^and_result116[200]^and_result116[201]^and_result116[202]^and_result116[203]^and_result116[204]^and_result116[205]^and_result116[206]^and_result116[207]^and_result116[208]^and_result116[209]^and_result116[210]^and_result116[211]^and_result116[212]^and_result116[213]^and_result116[214]^and_result116[215]^and_result116[216]^and_result116[217]^and_result116[218]^and_result116[219]^and_result116[220]^and_result116[221]^and_result116[222]^and_result116[223]^and_result116[224]^and_result116[225]^and_result116[226]^and_result116[227]^and_result116[228]^and_result116[229]^and_result116[230]^and_result116[231]^and_result116[232]^and_result116[233]^and_result116[234]^and_result116[235]^and_result116[236]^and_result116[237]^and_result116[238]^and_result116[239]^and_result116[240]^and_result116[241]^and_result116[242]^and_result116[243]^and_result116[244]^and_result116[245]^and_result116[246]^and_result116[247]^and_result116[248]^and_result116[249]^and_result116[250]^and_result116[251]^and_result116[252]^and_result116[253]^and_result116[254];
assign key[117]=and_result117[0]^and_result117[1]^and_result117[2]^and_result117[3]^and_result117[4]^and_result117[5]^and_result117[6]^and_result117[7]^and_result117[8]^and_result117[9]^and_result117[10]^and_result117[11]^and_result117[12]^and_result117[13]^and_result117[14]^and_result117[15]^and_result117[16]^and_result117[17]^and_result117[18]^and_result117[19]^and_result117[20]^and_result117[21]^and_result117[22]^and_result117[23]^and_result117[24]^and_result117[25]^and_result117[26]^and_result117[27]^and_result117[28]^and_result117[29]^and_result117[30]^and_result117[31]^and_result117[32]^and_result117[33]^and_result117[34]^and_result117[35]^and_result117[36]^and_result117[37]^and_result117[38]^and_result117[39]^and_result117[40]^and_result117[41]^and_result117[42]^and_result117[43]^and_result117[44]^and_result117[45]^and_result117[46]^and_result117[47]^and_result117[48]^and_result117[49]^and_result117[50]^and_result117[51]^and_result117[52]^and_result117[53]^and_result117[54]^and_result117[55]^and_result117[56]^and_result117[57]^and_result117[58]^and_result117[59]^and_result117[60]^and_result117[61]^and_result117[62]^and_result117[63]^and_result117[64]^and_result117[65]^and_result117[66]^and_result117[67]^and_result117[68]^and_result117[69]^and_result117[70]^and_result117[71]^and_result117[72]^and_result117[73]^and_result117[74]^and_result117[75]^and_result117[76]^and_result117[77]^and_result117[78]^and_result117[79]^and_result117[80]^and_result117[81]^and_result117[82]^and_result117[83]^and_result117[84]^and_result117[85]^and_result117[86]^and_result117[87]^and_result117[88]^and_result117[89]^and_result117[90]^and_result117[91]^and_result117[92]^and_result117[93]^and_result117[94]^and_result117[95]^and_result117[96]^and_result117[97]^and_result117[98]^and_result117[99]^and_result117[100]^and_result117[101]^and_result117[102]^and_result117[103]^and_result117[104]^and_result117[105]^and_result117[106]^and_result117[107]^and_result117[108]^and_result117[109]^and_result117[110]^and_result117[111]^and_result117[112]^and_result117[113]^and_result117[114]^and_result117[115]^and_result117[116]^and_result117[117]^and_result117[118]^and_result117[119]^and_result117[120]^and_result117[121]^and_result117[122]^and_result117[123]^and_result117[124]^and_result117[125]^and_result117[126]^and_result117[127]^and_result117[128]^and_result117[129]^and_result117[130]^and_result117[131]^and_result117[132]^and_result117[133]^and_result117[134]^and_result117[135]^and_result117[136]^and_result117[137]^and_result117[138]^and_result117[139]^and_result117[140]^and_result117[141]^and_result117[142]^and_result117[143]^and_result117[144]^and_result117[145]^and_result117[146]^and_result117[147]^and_result117[148]^and_result117[149]^and_result117[150]^and_result117[151]^and_result117[152]^and_result117[153]^and_result117[154]^and_result117[155]^and_result117[156]^and_result117[157]^and_result117[158]^and_result117[159]^and_result117[160]^and_result117[161]^and_result117[162]^and_result117[163]^and_result117[164]^and_result117[165]^and_result117[166]^and_result117[167]^and_result117[168]^and_result117[169]^and_result117[170]^and_result117[171]^and_result117[172]^and_result117[173]^and_result117[174]^and_result117[175]^and_result117[176]^and_result117[177]^and_result117[178]^and_result117[179]^and_result117[180]^and_result117[181]^and_result117[182]^and_result117[183]^and_result117[184]^and_result117[185]^and_result117[186]^and_result117[187]^and_result117[188]^and_result117[189]^and_result117[190]^and_result117[191]^and_result117[192]^and_result117[193]^and_result117[194]^and_result117[195]^and_result117[196]^and_result117[197]^and_result117[198]^and_result117[199]^and_result117[200]^and_result117[201]^and_result117[202]^and_result117[203]^and_result117[204]^and_result117[205]^and_result117[206]^and_result117[207]^and_result117[208]^and_result117[209]^and_result117[210]^and_result117[211]^and_result117[212]^and_result117[213]^and_result117[214]^and_result117[215]^and_result117[216]^and_result117[217]^and_result117[218]^and_result117[219]^and_result117[220]^and_result117[221]^and_result117[222]^and_result117[223]^and_result117[224]^and_result117[225]^and_result117[226]^and_result117[227]^and_result117[228]^and_result117[229]^and_result117[230]^and_result117[231]^and_result117[232]^and_result117[233]^and_result117[234]^and_result117[235]^and_result117[236]^and_result117[237]^and_result117[238]^and_result117[239]^and_result117[240]^and_result117[241]^and_result117[242]^and_result117[243]^and_result117[244]^and_result117[245]^and_result117[246]^and_result117[247]^and_result117[248]^and_result117[249]^and_result117[250]^and_result117[251]^and_result117[252]^and_result117[253]^and_result117[254];
assign key[118]=and_result118[0]^and_result118[1]^and_result118[2]^and_result118[3]^and_result118[4]^and_result118[5]^and_result118[6]^and_result118[7]^and_result118[8]^and_result118[9]^and_result118[10]^and_result118[11]^and_result118[12]^and_result118[13]^and_result118[14]^and_result118[15]^and_result118[16]^and_result118[17]^and_result118[18]^and_result118[19]^and_result118[20]^and_result118[21]^and_result118[22]^and_result118[23]^and_result118[24]^and_result118[25]^and_result118[26]^and_result118[27]^and_result118[28]^and_result118[29]^and_result118[30]^and_result118[31]^and_result118[32]^and_result118[33]^and_result118[34]^and_result118[35]^and_result118[36]^and_result118[37]^and_result118[38]^and_result118[39]^and_result118[40]^and_result118[41]^and_result118[42]^and_result118[43]^and_result118[44]^and_result118[45]^and_result118[46]^and_result118[47]^and_result118[48]^and_result118[49]^and_result118[50]^and_result118[51]^and_result118[52]^and_result118[53]^and_result118[54]^and_result118[55]^and_result118[56]^and_result118[57]^and_result118[58]^and_result118[59]^and_result118[60]^and_result118[61]^and_result118[62]^and_result118[63]^and_result118[64]^and_result118[65]^and_result118[66]^and_result118[67]^and_result118[68]^and_result118[69]^and_result118[70]^and_result118[71]^and_result118[72]^and_result118[73]^and_result118[74]^and_result118[75]^and_result118[76]^and_result118[77]^and_result118[78]^and_result118[79]^and_result118[80]^and_result118[81]^and_result118[82]^and_result118[83]^and_result118[84]^and_result118[85]^and_result118[86]^and_result118[87]^and_result118[88]^and_result118[89]^and_result118[90]^and_result118[91]^and_result118[92]^and_result118[93]^and_result118[94]^and_result118[95]^and_result118[96]^and_result118[97]^and_result118[98]^and_result118[99]^and_result118[100]^and_result118[101]^and_result118[102]^and_result118[103]^and_result118[104]^and_result118[105]^and_result118[106]^and_result118[107]^and_result118[108]^and_result118[109]^and_result118[110]^and_result118[111]^and_result118[112]^and_result118[113]^and_result118[114]^and_result118[115]^and_result118[116]^and_result118[117]^and_result118[118]^and_result118[119]^and_result118[120]^and_result118[121]^and_result118[122]^and_result118[123]^and_result118[124]^and_result118[125]^and_result118[126]^and_result118[127]^and_result118[128]^and_result118[129]^and_result118[130]^and_result118[131]^and_result118[132]^and_result118[133]^and_result118[134]^and_result118[135]^and_result118[136]^and_result118[137]^and_result118[138]^and_result118[139]^and_result118[140]^and_result118[141]^and_result118[142]^and_result118[143]^and_result118[144]^and_result118[145]^and_result118[146]^and_result118[147]^and_result118[148]^and_result118[149]^and_result118[150]^and_result118[151]^and_result118[152]^and_result118[153]^and_result118[154]^and_result118[155]^and_result118[156]^and_result118[157]^and_result118[158]^and_result118[159]^and_result118[160]^and_result118[161]^and_result118[162]^and_result118[163]^and_result118[164]^and_result118[165]^and_result118[166]^and_result118[167]^and_result118[168]^and_result118[169]^and_result118[170]^and_result118[171]^and_result118[172]^and_result118[173]^and_result118[174]^and_result118[175]^and_result118[176]^and_result118[177]^and_result118[178]^and_result118[179]^and_result118[180]^and_result118[181]^and_result118[182]^and_result118[183]^and_result118[184]^and_result118[185]^and_result118[186]^and_result118[187]^and_result118[188]^and_result118[189]^and_result118[190]^and_result118[191]^and_result118[192]^and_result118[193]^and_result118[194]^and_result118[195]^and_result118[196]^and_result118[197]^and_result118[198]^and_result118[199]^and_result118[200]^and_result118[201]^and_result118[202]^and_result118[203]^and_result118[204]^and_result118[205]^and_result118[206]^and_result118[207]^and_result118[208]^and_result118[209]^and_result118[210]^and_result118[211]^and_result118[212]^and_result118[213]^and_result118[214]^and_result118[215]^and_result118[216]^and_result118[217]^and_result118[218]^and_result118[219]^and_result118[220]^and_result118[221]^and_result118[222]^and_result118[223]^and_result118[224]^and_result118[225]^and_result118[226]^and_result118[227]^and_result118[228]^and_result118[229]^and_result118[230]^and_result118[231]^and_result118[232]^and_result118[233]^and_result118[234]^and_result118[235]^and_result118[236]^and_result118[237]^and_result118[238]^and_result118[239]^and_result118[240]^and_result118[241]^and_result118[242]^and_result118[243]^and_result118[244]^and_result118[245]^and_result118[246]^and_result118[247]^and_result118[248]^and_result118[249]^and_result118[250]^and_result118[251]^and_result118[252]^and_result118[253]^and_result118[254];
assign key[119]=and_result119[0]^and_result119[1]^and_result119[2]^and_result119[3]^and_result119[4]^and_result119[5]^and_result119[6]^and_result119[7]^and_result119[8]^and_result119[9]^and_result119[10]^and_result119[11]^and_result119[12]^and_result119[13]^and_result119[14]^and_result119[15]^and_result119[16]^and_result119[17]^and_result119[18]^and_result119[19]^and_result119[20]^and_result119[21]^and_result119[22]^and_result119[23]^and_result119[24]^and_result119[25]^and_result119[26]^and_result119[27]^and_result119[28]^and_result119[29]^and_result119[30]^and_result119[31]^and_result119[32]^and_result119[33]^and_result119[34]^and_result119[35]^and_result119[36]^and_result119[37]^and_result119[38]^and_result119[39]^and_result119[40]^and_result119[41]^and_result119[42]^and_result119[43]^and_result119[44]^and_result119[45]^and_result119[46]^and_result119[47]^and_result119[48]^and_result119[49]^and_result119[50]^and_result119[51]^and_result119[52]^and_result119[53]^and_result119[54]^and_result119[55]^and_result119[56]^and_result119[57]^and_result119[58]^and_result119[59]^and_result119[60]^and_result119[61]^and_result119[62]^and_result119[63]^and_result119[64]^and_result119[65]^and_result119[66]^and_result119[67]^and_result119[68]^and_result119[69]^and_result119[70]^and_result119[71]^and_result119[72]^and_result119[73]^and_result119[74]^and_result119[75]^and_result119[76]^and_result119[77]^and_result119[78]^and_result119[79]^and_result119[80]^and_result119[81]^and_result119[82]^and_result119[83]^and_result119[84]^and_result119[85]^and_result119[86]^and_result119[87]^and_result119[88]^and_result119[89]^and_result119[90]^and_result119[91]^and_result119[92]^and_result119[93]^and_result119[94]^and_result119[95]^and_result119[96]^and_result119[97]^and_result119[98]^and_result119[99]^and_result119[100]^and_result119[101]^and_result119[102]^and_result119[103]^and_result119[104]^and_result119[105]^and_result119[106]^and_result119[107]^and_result119[108]^and_result119[109]^and_result119[110]^and_result119[111]^and_result119[112]^and_result119[113]^and_result119[114]^and_result119[115]^and_result119[116]^and_result119[117]^and_result119[118]^and_result119[119]^and_result119[120]^and_result119[121]^and_result119[122]^and_result119[123]^and_result119[124]^and_result119[125]^and_result119[126]^and_result119[127]^and_result119[128]^and_result119[129]^and_result119[130]^and_result119[131]^and_result119[132]^and_result119[133]^and_result119[134]^and_result119[135]^and_result119[136]^and_result119[137]^and_result119[138]^and_result119[139]^and_result119[140]^and_result119[141]^and_result119[142]^and_result119[143]^and_result119[144]^and_result119[145]^and_result119[146]^and_result119[147]^and_result119[148]^and_result119[149]^and_result119[150]^and_result119[151]^and_result119[152]^and_result119[153]^and_result119[154]^and_result119[155]^and_result119[156]^and_result119[157]^and_result119[158]^and_result119[159]^and_result119[160]^and_result119[161]^and_result119[162]^and_result119[163]^and_result119[164]^and_result119[165]^and_result119[166]^and_result119[167]^and_result119[168]^and_result119[169]^and_result119[170]^and_result119[171]^and_result119[172]^and_result119[173]^and_result119[174]^and_result119[175]^and_result119[176]^and_result119[177]^and_result119[178]^and_result119[179]^and_result119[180]^and_result119[181]^and_result119[182]^and_result119[183]^and_result119[184]^and_result119[185]^and_result119[186]^and_result119[187]^and_result119[188]^and_result119[189]^and_result119[190]^and_result119[191]^and_result119[192]^and_result119[193]^and_result119[194]^and_result119[195]^and_result119[196]^and_result119[197]^and_result119[198]^and_result119[199]^and_result119[200]^and_result119[201]^and_result119[202]^and_result119[203]^and_result119[204]^and_result119[205]^and_result119[206]^and_result119[207]^and_result119[208]^and_result119[209]^and_result119[210]^and_result119[211]^and_result119[212]^and_result119[213]^and_result119[214]^and_result119[215]^and_result119[216]^and_result119[217]^and_result119[218]^and_result119[219]^and_result119[220]^and_result119[221]^and_result119[222]^and_result119[223]^and_result119[224]^and_result119[225]^and_result119[226]^and_result119[227]^and_result119[228]^and_result119[229]^and_result119[230]^and_result119[231]^and_result119[232]^and_result119[233]^and_result119[234]^and_result119[235]^and_result119[236]^and_result119[237]^and_result119[238]^and_result119[239]^and_result119[240]^and_result119[241]^and_result119[242]^and_result119[243]^and_result119[244]^and_result119[245]^and_result119[246]^and_result119[247]^and_result119[248]^and_result119[249]^and_result119[250]^and_result119[251]^and_result119[252]^and_result119[253]^and_result119[254];
assign key[120]=and_result120[0]^and_result120[1]^and_result120[2]^and_result120[3]^and_result120[4]^and_result120[5]^and_result120[6]^and_result120[7]^and_result120[8]^and_result120[9]^and_result120[10]^and_result120[11]^and_result120[12]^and_result120[13]^and_result120[14]^and_result120[15]^and_result120[16]^and_result120[17]^and_result120[18]^and_result120[19]^and_result120[20]^and_result120[21]^and_result120[22]^and_result120[23]^and_result120[24]^and_result120[25]^and_result120[26]^and_result120[27]^and_result120[28]^and_result120[29]^and_result120[30]^and_result120[31]^and_result120[32]^and_result120[33]^and_result120[34]^and_result120[35]^and_result120[36]^and_result120[37]^and_result120[38]^and_result120[39]^and_result120[40]^and_result120[41]^and_result120[42]^and_result120[43]^and_result120[44]^and_result120[45]^and_result120[46]^and_result120[47]^and_result120[48]^and_result120[49]^and_result120[50]^and_result120[51]^and_result120[52]^and_result120[53]^and_result120[54]^and_result120[55]^and_result120[56]^and_result120[57]^and_result120[58]^and_result120[59]^and_result120[60]^and_result120[61]^and_result120[62]^and_result120[63]^and_result120[64]^and_result120[65]^and_result120[66]^and_result120[67]^and_result120[68]^and_result120[69]^and_result120[70]^and_result120[71]^and_result120[72]^and_result120[73]^and_result120[74]^and_result120[75]^and_result120[76]^and_result120[77]^and_result120[78]^and_result120[79]^and_result120[80]^and_result120[81]^and_result120[82]^and_result120[83]^and_result120[84]^and_result120[85]^and_result120[86]^and_result120[87]^and_result120[88]^and_result120[89]^and_result120[90]^and_result120[91]^and_result120[92]^and_result120[93]^and_result120[94]^and_result120[95]^and_result120[96]^and_result120[97]^and_result120[98]^and_result120[99]^and_result120[100]^and_result120[101]^and_result120[102]^and_result120[103]^and_result120[104]^and_result120[105]^and_result120[106]^and_result120[107]^and_result120[108]^and_result120[109]^and_result120[110]^and_result120[111]^and_result120[112]^and_result120[113]^and_result120[114]^and_result120[115]^and_result120[116]^and_result120[117]^and_result120[118]^and_result120[119]^and_result120[120]^and_result120[121]^and_result120[122]^and_result120[123]^and_result120[124]^and_result120[125]^and_result120[126]^and_result120[127]^and_result120[128]^and_result120[129]^and_result120[130]^and_result120[131]^and_result120[132]^and_result120[133]^and_result120[134]^and_result120[135]^and_result120[136]^and_result120[137]^and_result120[138]^and_result120[139]^and_result120[140]^and_result120[141]^and_result120[142]^and_result120[143]^and_result120[144]^and_result120[145]^and_result120[146]^and_result120[147]^and_result120[148]^and_result120[149]^and_result120[150]^and_result120[151]^and_result120[152]^and_result120[153]^and_result120[154]^and_result120[155]^and_result120[156]^and_result120[157]^and_result120[158]^and_result120[159]^and_result120[160]^and_result120[161]^and_result120[162]^and_result120[163]^and_result120[164]^and_result120[165]^and_result120[166]^and_result120[167]^and_result120[168]^and_result120[169]^and_result120[170]^and_result120[171]^and_result120[172]^and_result120[173]^and_result120[174]^and_result120[175]^and_result120[176]^and_result120[177]^and_result120[178]^and_result120[179]^and_result120[180]^and_result120[181]^and_result120[182]^and_result120[183]^and_result120[184]^and_result120[185]^and_result120[186]^and_result120[187]^and_result120[188]^and_result120[189]^and_result120[190]^and_result120[191]^and_result120[192]^and_result120[193]^and_result120[194]^and_result120[195]^and_result120[196]^and_result120[197]^and_result120[198]^and_result120[199]^and_result120[200]^and_result120[201]^and_result120[202]^and_result120[203]^and_result120[204]^and_result120[205]^and_result120[206]^and_result120[207]^and_result120[208]^and_result120[209]^and_result120[210]^and_result120[211]^and_result120[212]^and_result120[213]^and_result120[214]^and_result120[215]^and_result120[216]^and_result120[217]^and_result120[218]^and_result120[219]^and_result120[220]^and_result120[221]^and_result120[222]^and_result120[223]^and_result120[224]^and_result120[225]^and_result120[226]^and_result120[227]^and_result120[228]^and_result120[229]^and_result120[230]^and_result120[231]^and_result120[232]^and_result120[233]^and_result120[234]^and_result120[235]^and_result120[236]^and_result120[237]^and_result120[238]^and_result120[239]^and_result120[240]^and_result120[241]^and_result120[242]^and_result120[243]^and_result120[244]^and_result120[245]^and_result120[246]^and_result120[247]^and_result120[248]^and_result120[249]^and_result120[250]^and_result120[251]^and_result120[252]^and_result120[253]^and_result120[254];
assign key[121]=and_result121[0]^and_result121[1]^and_result121[2]^and_result121[3]^and_result121[4]^and_result121[5]^and_result121[6]^and_result121[7]^and_result121[8]^and_result121[9]^and_result121[10]^and_result121[11]^and_result121[12]^and_result121[13]^and_result121[14]^and_result121[15]^and_result121[16]^and_result121[17]^and_result121[18]^and_result121[19]^and_result121[20]^and_result121[21]^and_result121[22]^and_result121[23]^and_result121[24]^and_result121[25]^and_result121[26]^and_result121[27]^and_result121[28]^and_result121[29]^and_result121[30]^and_result121[31]^and_result121[32]^and_result121[33]^and_result121[34]^and_result121[35]^and_result121[36]^and_result121[37]^and_result121[38]^and_result121[39]^and_result121[40]^and_result121[41]^and_result121[42]^and_result121[43]^and_result121[44]^and_result121[45]^and_result121[46]^and_result121[47]^and_result121[48]^and_result121[49]^and_result121[50]^and_result121[51]^and_result121[52]^and_result121[53]^and_result121[54]^and_result121[55]^and_result121[56]^and_result121[57]^and_result121[58]^and_result121[59]^and_result121[60]^and_result121[61]^and_result121[62]^and_result121[63]^and_result121[64]^and_result121[65]^and_result121[66]^and_result121[67]^and_result121[68]^and_result121[69]^and_result121[70]^and_result121[71]^and_result121[72]^and_result121[73]^and_result121[74]^and_result121[75]^and_result121[76]^and_result121[77]^and_result121[78]^and_result121[79]^and_result121[80]^and_result121[81]^and_result121[82]^and_result121[83]^and_result121[84]^and_result121[85]^and_result121[86]^and_result121[87]^and_result121[88]^and_result121[89]^and_result121[90]^and_result121[91]^and_result121[92]^and_result121[93]^and_result121[94]^and_result121[95]^and_result121[96]^and_result121[97]^and_result121[98]^and_result121[99]^and_result121[100]^and_result121[101]^and_result121[102]^and_result121[103]^and_result121[104]^and_result121[105]^and_result121[106]^and_result121[107]^and_result121[108]^and_result121[109]^and_result121[110]^and_result121[111]^and_result121[112]^and_result121[113]^and_result121[114]^and_result121[115]^and_result121[116]^and_result121[117]^and_result121[118]^and_result121[119]^and_result121[120]^and_result121[121]^and_result121[122]^and_result121[123]^and_result121[124]^and_result121[125]^and_result121[126]^and_result121[127]^and_result121[128]^and_result121[129]^and_result121[130]^and_result121[131]^and_result121[132]^and_result121[133]^and_result121[134]^and_result121[135]^and_result121[136]^and_result121[137]^and_result121[138]^and_result121[139]^and_result121[140]^and_result121[141]^and_result121[142]^and_result121[143]^and_result121[144]^and_result121[145]^and_result121[146]^and_result121[147]^and_result121[148]^and_result121[149]^and_result121[150]^and_result121[151]^and_result121[152]^and_result121[153]^and_result121[154]^and_result121[155]^and_result121[156]^and_result121[157]^and_result121[158]^and_result121[159]^and_result121[160]^and_result121[161]^and_result121[162]^and_result121[163]^and_result121[164]^and_result121[165]^and_result121[166]^and_result121[167]^and_result121[168]^and_result121[169]^and_result121[170]^and_result121[171]^and_result121[172]^and_result121[173]^and_result121[174]^and_result121[175]^and_result121[176]^and_result121[177]^and_result121[178]^and_result121[179]^and_result121[180]^and_result121[181]^and_result121[182]^and_result121[183]^and_result121[184]^and_result121[185]^and_result121[186]^and_result121[187]^and_result121[188]^and_result121[189]^and_result121[190]^and_result121[191]^and_result121[192]^and_result121[193]^and_result121[194]^and_result121[195]^and_result121[196]^and_result121[197]^and_result121[198]^and_result121[199]^and_result121[200]^and_result121[201]^and_result121[202]^and_result121[203]^and_result121[204]^and_result121[205]^and_result121[206]^and_result121[207]^and_result121[208]^and_result121[209]^and_result121[210]^and_result121[211]^and_result121[212]^and_result121[213]^and_result121[214]^and_result121[215]^and_result121[216]^and_result121[217]^and_result121[218]^and_result121[219]^and_result121[220]^and_result121[221]^and_result121[222]^and_result121[223]^and_result121[224]^and_result121[225]^and_result121[226]^and_result121[227]^and_result121[228]^and_result121[229]^and_result121[230]^and_result121[231]^and_result121[232]^and_result121[233]^and_result121[234]^and_result121[235]^and_result121[236]^and_result121[237]^and_result121[238]^and_result121[239]^and_result121[240]^and_result121[241]^and_result121[242]^and_result121[243]^and_result121[244]^and_result121[245]^and_result121[246]^and_result121[247]^and_result121[248]^and_result121[249]^and_result121[250]^and_result121[251]^and_result121[252]^and_result121[253]^and_result121[254];
assign key[122]=and_result122[0]^and_result122[1]^and_result122[2]^and_result122[3]^and_result122[4]^and_result122[5]^and_result122[6]^and_result122[7]^and_result122[8]^and_result122[9]^and_result122[10]^and_result122[11]^and_result122[12]^and_result122[13]^and_result122[14]^and_result122[15]^and_result122[16]^and_result122[17]^and_result122[18]^and_result122[19]^and_result122[20]^and_result122[21]^and_result122[22]^and_result122[23]^and_result122[24]^and_result122[25]^and_result122[26]^and_result122[27]^and_result122[28]^and_result122[29]^and_result122[30]^and_result122[31]^and_result122[32]^and_result122[33]^and_result122[34]^and_result122[35]^and_result122[36]^and_result122[37]^and_result122[38]^and_result122[39]^and_result122[40]^and_result122[41]^and_result122[42]^and_result122[43]^and_result122[44]^and_result122[45]^and_result122[46]^and_result122[47]^and_result122[48]^and_result122[49]^and_result122[50]^and_result122[51]^and_result122[52]^and_result122[53]^and_result122[54]^and_result122[55]^and_result122[56]^and_result122[57]^and_result122[58]^and_result122[59]^and_result122[60]^and_result122[61]^and_result122[62]^and_result122[63]^and_result122[64]^and_result122[65]^and_result122[66]^and_result122[67]^and_result122[68]^and_result122[69]^and_result122[70]^and_result122[71]^and_result122[72]^and_result122[73]^and_result122[74]^and_result122[75]^and_result122[76]^and_result122[77]^and_result122[78]^and_result122[79]^and_result122[80]^and_result122[81]^and_result122[82]^and_result122[83]^and_result122[84]^and_result122[85]^and_result122[86]^and_result122[87]^and_result122[88]^and_result122[89]^and_result122[90]^and_result122[91]^and_result122[92]^and_result122[93]^and_result122[94]^and_result122[95]^and_result122[96]^and_result122[97]^and_result122[98]^and_result122[99]^and_result122[100]^and_result122[101]^and_result122[102]^and_result122[103]^and_result122[104]^and_result122[105]^and_result122[106]^and_result122[107]^and_result122[108]^and_result122[109]^and_result122[110]^and_result122[111]^and_result122[112]^and_result122[113]^and_result122[114]^and_result122[115]^and_result122[116]^and_result122[117]^and_result122[118]^and_result122[119]^and_result122[120]^and_result122[121]^and_result122[122]^and_result122[123]^and_result122[124]^and_result122[125]^and_result122[126]^and_result122[127]^and_result122[128]^and_result122[129]^and_result122[130]^and_result122[131]^and_result122[132]^and_result122[133]^and_result122[134]^and_result122[135]^and_result122[136]^and_result122[137]^and_result122[138]^and_result122[139]^and_result122[140]^and_result122[141]^and_result122[142]^and_result122[143]^and_result122[144]^and_result122[145]^and_result122[146]^and_result122[147]^and_result122[148]^and_result122[149]^and_result122[150]^and_result122[151]^and_result122[152]^and_result122[153]^and_result122[154]^and_result122[155]^and_result122[156]^and_result122[157]^and_result122[158]^and_result122[159]^and_result122[160]^and_result122[161]^and_result122[162]^and_result122[163]^and_result122[164]^and_result122[165]^and_result122[166]^and_result122[167]^and_result122[168]^and_result122[169]^and_result122[170]^and_result122[171]^and_result122[172]^and_result122[173]^and_result122[174]^and_result122[175]^and_result122[176]^and_result122[177]^and_result122[178]^and_result122[179]^and_result122[180]^and_result122[181]^and_result122[182]^and_result122[183]^and_result122[184]^and_result122[185]^and_result122[186]^and_result122[187]^and_result122[188]^and_result122[189]^and_result122[190]^and_result122[191]^and_result122[192]^and_result122[193]^and_result122[194]^and_result122[195]^and_result122[196]^and_result122[197]^and_result122[198]^and_result122[199]^and_result122[200]^and_result122[201]^and_result122[202]^and_result122[203]^and_result122[204]^and_result122[205]^and_result122[206]^and_result122[207]^and_result122[208]^and_result122[209]^and_result122[210]^and_result122[211]^and_result122[212]^and_result122[213]^and_result122[214]^and_result122[215]^and_result122[216]^and_result122[217]^and_result122[218]^and_result122[219]^and_result122[220]^and_result122[221]^and_result122[222]^and_result122[223]^and_result122[224]^and_result122[225]^and_result122[226]^and_result122[227]^and_result122[228]^and_result122[229]^and_result122[230]^and_result122[231]^and_result122[232]^and_result122[233]^and_result122[234]^and_result122[235]^and_result122[236]^and_result122[237]^and_result122[238]^and_result122[239]^and_result122[240]^and_result122[241]^and_result122[242]^and_result122[243]^and_result122[244]^and_result122[245]^and_result122[246]^and_result122[247]^and_result122[248]^and_result122[249]^and_result122[250]^and_result122[251]^and_result122[252]^and_result122[253]^and_result122[254];
assign key[123]=and_result123[0]^and_result123[1]^and_result123[2]^and_result123[3]^and_result123[4]^and_result123[5]^and_result123[6]^and_result123[7]^and_result123[8]^and_result123[9]^and_result123[10]^and_result123[11]^and_result123[12]^and_result123[13]^and_result123[14]^and_result123[15]^and_result123[16]^and_result123[17]^and_result123[18]^and_result123[19]^and_result123[20]^and_result123[21]^and_result123[22]^and_result123[23]^and_result123[24]^and_result123[25]^and_result123[26]^and_result123[27]^and_result123[28]^and_result123[29]^and_result123[30]^and_result123[31]^and_result123[32]^and_result123[33]^and_result123[34]^and_result123[35]^and_result123[36]^and_result123[37]^and_result123[38]^and_result123[39]^and_result123[40]^and_result123[41]^and_result123[42]^and_result123[43]^and_result123[44]^and_result123[45]^and_result123[46]^and_result123[47]^and_result123[48]^and_result123[49]^and_result123[50]^and_result123[51]^and_result123[52]^and_result123[53]^and_result123[54]^and_result123[55]^and_result123[56]^and_result123[57]^and_result123[58]^and_result123[59]^and_result123[60]^and_result123[61]^and_result123[62]^and_result123[63]^and_result123[64]^and_result123[65]^and_result123[66]^and_result123[67]^and_result123[68]^and_result123[69]^and_result123[70]^and_result123[71]^and_result123[72]^and_result123[73]^and_result123[74]^and_result123[75]^and_result123[76]^and_result123[77]^and_result123[78]^and_result123[79]^and_result123[80]^and_result123[81]^and_result123[82]^and_result123[83]^and_result123[84]^and_result123[85]^and_result123[86]^and_result123[87]^and_result123[88]^and_result123[89]^and_result123[90]^and_result123[91]^and_result123[92]^and_result123[93]^and_result123[94]^and_result123[95]^and_result123[96]^and_result123[97]^and_result123[98]^and_result123[99]^and_result123[100]^and_result123[101]^and_result123[102]^and_result123[103]^and_result123[104]^and_result123[105]^and_result123[106]^and_result123[107]^and_result123[108]^and_result123[109]^and_result123[110]^and_result123[111]^and_result123[112]^and_result123[113]^and_result123[114]^and_result123[115]^and_result123[116]^and_result123[117]^and_result123[118]^and_result123[119]^and_result123[120]^and_result123[121]^and_result123[122]^and_result123[123]^and_result123[124]^and_result123[125]^and_result123[126]^and_result123[127]^and_result123[128]^and_result123[129]^and_result123[130]^and_result123[131]^and_result123[132]^and_result123[133]^and_result123[134]^and_result123[135]^and_result123[136]^and_result123[137]^and_result123[138]^and_result123[139]^and_result123[140]^and_result123[141]^and_result123[142]^and_result123[143]^and_result123[144]^and_result123[145]^and_result123[146]^and_result123[147]^and_result123[148]^and_result123[149]^and_result123[150]^and_result123[151]^and_result123[152]^and_result123[153]^and_result123[154]^and_result123[155]^and_result123[156]^and_result123[157]^and_result123[158]^and_result123[159]^and_result123[160]^and_result123[161]^and_result123[162]^and_result123[163]^and_result123[164]^and_result123[165]^and_result123[166]^and_result123[167]^and_result123[168]^and_result123[169]^and_result123[170]^and_result123[171]^and_result123[172]^and_result123[173]^and_result123[174]^and_result123[175]^and_result123[176]^and_result123[177]^and_result123[178]^and_result123[179]^and_result123[180]^and_result123[181]^and_result123[182]^and_result123[183]^and_result123[184]^and_result123[185]^and_result123[186]^and_result123[187]^and_result123[188]^and_result123[189]^and_result123[190]^and_result123[191]^and_result123[192]^and_result123[193]^and_result123[194]^and_result123[195]^and_result123[196]^and_result123[197]^and_result123[198]^and_result123[199]^and_result123[200]^and_result123[201]^and_result123[202]^and_result123[203]^and_result123[204]^and_result123[205]^and_result123[206]^and_result123[207]^and_result123[208]^and_result123[209]^and_result123[210]^and_result123[211]^and_result123[212]^and_result123[213]^and_result123[214]^and_result123[215]^and_result123[216]^and_result123[217]^and_result123[218]^and_result123[219]^and_result123[220]^and_result123[221]^and_result123[222]^and_result123[223]^and_result123[224]^and_result123[225]^and_result123[226]^and_result123[227]^and_result123[228]^and_result123[229]^and_result123[230]^and_result123[231]^and_result123[232]^and_result123[233]^and_result123[234]^and_result123[235]^and_result123[236]^and_result123[237]^and_result123[238]^and_result123[239]^and_result123[240]^and_result123[241]^and_result123[242]^and_result123[243]^and_result123[244]^and_result123[245]^and_result123[246]^and_result123[247]^and_result123[248]^and_result123[249]^and_result123[250]^and_result123[251]^and_result123[252]^and_result123[253]^and_result123[254];
assign key[124]=and_result124[0]^and_result124[1]^and_result124[2]^and_result124[3]^and_result124[4]^and_result124[5]^and_result124[6]^and_result124[7]^and_result124[8]^and_result124[9]^and_result124[10]^and_result124[11]^and_result124[12]^and_result124[13]^and_result124[14]^and_result124[15]^and_result124[16]^and_result124[17]^and_result124[18]^and_result124[19]^and_result124[20]^and_result124[21]^and_result124[22]^and_result124[23]^and_result124[24]^and_result124[25]^and_result124[26]^and_result124[27]^and_result124[28]^and_result124[29]^and_result124[30]^and_result124[31]^and_result124[32]^and_result124[33]^and_result124[34]^and_result124[35]^and_result124[36]^and_result124[37]^and_result124[38]^and_result124[39]^and_result124[40]^and_result124[41]^and_result124[42]^and_result124[43]^and_result124[44]^and_result124[45]^and_result124[46]^and_result124[47]^and_result124[48]^and_result124[49]^and_result124[50]^and_result124[51]^and_result124[52]^and_result124[53]^and_result124[54]^and_result124[55]^and_result124[56]^and_result124[57]^and_result124[58]^and_result124[59]^and_result124[60]^and_result124[61]^and_result124[62]^and_result124[63]^and_result124[64]^and_result124[65]^and_result124[66]^and_result124[67]^and_result124[68]^and_result124[69]^and_result124[70]^and_result124[71]^and_result124[72]^and_result124[73]^and_result124[74]^and_result124[75]^and_result124[76]^and_result124[77]^and_result124[78]^and_result124[79]^and_result124[80]^and_result124[81]^and_result124[82]^and_result124[83]^and_result124[84]^and_result124[85]^and_result124[86]^and_result124[87]^and_result124[88]^and_result124[89]^and_result124[90]^and_result124[91]^and_result124[92]^and_result124[93]^and_result124[94]^and_result124[95]^and_result124[96]^and_result124[97]^and_result124[98]^and_result124[99]^and_result124[100]^and_result124[101]^and_result124[102]^and_result124[103]^and_result124[104]^and_result124[105]^and_result124[106]^and_result124[107]^and_result124[108]^and_result124[109]^and_result124[110]^and_result124[111]^and_result124[112]^and_result124[113]^and_result124[114]^and_result124[115]^and_result124[116]^and_result124[117]^and_result124[118]^and_result124[119]^and_result124[120]^and_result124[121]^and_result124[122]^and_result124[123]^and_result124[124]^and_result124[125]^and_result124[126]^and_result124[127]^and_result124[128]^and_result124[129]^and_result124[130]^and_result124[131]^and_result124[132]^and_result124[133]^and_result124[134]^and_result124[135]^and_result124[136]^and_result124[137]^and_result124[138]^and_result124[139]^and_result124[140]^and_result124[141]^and_result124[142]^and_result124[143]^and_result124[144]^and_result124[145]^and_result124[146]^and_result124[147]^and_result124[148]^and_result124[149]^and_result124[150]^and_result124[151]^and_result124[152]^and_result124[153]^and_result124[154]^and_result124[155]^and_result124[156]^and_result124[157]^and_result124[158]^and_result124[159]^and_result124[160]^and_result124[161]^and_result124[162]^and_result124[163]^and_result124[164]^and_result124[165]^and_result124[166]^and_result124[167]^and_result124[168]^and_result124[169]^and_result124[170]^and_result124[171]^and_result124[172]^and_result124[173]^and_result124[174]^and_result124[175]^and_result124[176]^and_result124[177]^and_result124[178]^and_result124[179]^and_result124[180]^and_result124[181]^and_result124[182]^and_result124[183]^and_result124[184]^and_result124[185]^and_result124[186]^and_result124[187]^and_result124[188]^and_result124[189]^and_result124[190]^and_result124[191]^and_result124[192]^and_result124[193]^and_result124[194]^and_result124[195]^and_result124[196]^and_result124[197]^and_result124[198]^and_result124[199]^and_result124[200]^and_result124[201]^and_result124[202]^and_result124[203]^and_result124[204]^and_result124[205]^and_result124[206]^and_result124[207]^and_result124[208]^and_result124[209]^and_result124[210]^and_result124[211]^and_result124[212]^and_result124[213]^and_result124[214]^and_result124[215]^and_result124[216]^and_result124[217]^and_result124[218]^and_result124[219]^and_result124[220]^and_result124[221]^and_result124[222]^and_result124[223]^and_result124[224]^and_result124[225]^and_result124[226]^and_result124[227]^and_result124[228]^and_result124[229]^and_result124[230]^and_result124[231]^and_result124[232]^and_result124[233]^and_result124[234]^and_result124[235]^and_result124[236]^and_result124[237]^and_result124[238]^and_result124[239]^and_result124[240]^and_result124[241]^and_result124[242]^and_result124[243]^and_result124[244]^and_result124[245]^and_result124[246]^and_result124[247]^and_result124[248]^and_result124[249]^and_result124[250]^and_result124[251]^and_result124[252]^and_result124[253]^and_result124[254];
assign key[125]=and_result125[0]^and_result125[1]^and_result125[2]^and_result125[3]^and_result125[4]^and_result125[5]^and_result125[6]^and_result125[7]^and_result125[8]^and_result125[9]^and_result125[10]^and_result125[11]^and_result125[12]^and_result125[13]^and_result125[14]^and_result125[15]^and_result125[16]^and_result125[17]^and_result125[18]^and_result125[19]^and_result125[20]^and_result125[21]^and_result125[22]^and_result125[23]^and_result125[24]^and_result125[25]^and_result125[26]^and_result125[27]^and_result125[28]^and_result125[29]^and_result125[30]^and_result125[31]^and_result125[32]^and_result125[33]^and_result125[34]^and_result125[35]^and_result125[36]^and_result125[37]^and_result125[38]^and_result125[39]^and_result125[40]^and_result125[41]^and_result125[42]^and_result125[43]^and_result125[44]^and_result125[45]^and_result125[46]^and_result125[47]^and_result125[48]^and_result125[49]^and_result125[50]^and_result125[51]^and_result125[52]^and_result125[53]^and_result125[54]^and_result125[55]^and_result125[56]^and_result125[57]^and_result125[58]^and_result125[59]^and_result125[60]^and_result125[61]^and_result125[62]^and_result125[63]^and_result125[64]^and_result125[65]^and_result125[66]^and_result125[67]^and_result125[68]^and_result125[69]^and_result125[70]^and_result125[71]^and_result125[72]^and_result125[73]^and_result125[74]^and_result125[75]^and_result125[76]^and_result125[77]^and_result125[78]^and_result125[79]^and_result125[80]^and_result125[81]^and_result125[82]^and_result125[83]^and_result125[84]^and_result125[85]^and_result125[86]^and_result125[87]^and_result125[88]^and_result125[89]^and_result125[90]^and_result125[91]^and_result125[92]^and_result125[93]^and_result125[94]^and_result125[95]^and_result125[96]^and_result125[97]^and_result125[98]^and_result125[99]^and_result125[100]^and_result125[101]^and_result125[102]^and_result125[103]^and_result125[104]^and_result125[105]^and_result125[106]^and_result125[107]^and_result125[108]^and_result125[109]^and_result125[110]^and_result125[111]^and_result125[112]^and_result125[113]^and_result125[114]^and_result125[115]^and_result125[116]^and_result125[117]^and_result125[118]^and_result125[119]^and_result125[120]^and_result125[121]^and_result125[122]^and_result125[123]^and_result125[124]^and_result125[125]^and_result125[126]^and_result125[127]^and_result125[128]^and_result125[129]^and_result125[130]^and_result125[131]^and_result125[132]^and_result125[133]^and_result125[134]^and_result125[135]^and_result125[136]^and_result125[137]^and_result125[138]^and_result125[139]^and_result125[140]^and_result125[141]^and_result125[142]^and_result125[143]^and_result125[144]^and_result125[145]^and_result125[146]^and_result125[147]^and_result125[148]^and_result125[149]^and_result125[150]^and_result125[151]^and_result125[152]^and_result125[153]^and_result125[154]^and_result125[155]^and_result125[156]^and_result125[157]^and_result125[158]^and_result125[159]^and_result125[160]^and_result125[161]^and_result125[162]^and_result125[163]^and_result125[164]^and_result125[165]^and_result125[166]^and_result125[167]^and_result125[168]^and_result125[169]^and_result125[170]^and_result125[171]^and_result125[172]^and_result125[173]^and_result125[174]^and_result125[175]^and_result125[176]^and_result125[177]^and_result125[178]^and_result125[179]^and_result125[180]^and_result125[181]^and_result125[182]^and_result125[183]^and_result125[184]^and_result125[185]^and_result125[186]^and_result125[187]^and_result125[188]^and_result125[189]^and_result125[190]^and_result125[191]^and_result125[192]^and_result125[193]^and_result125[194]^and_result125[195]^and_result125[196]^and_result125[197]^and_result125[198]^and_result125[199]^and_result125[200]^and_result125[201]^and_result125[202]^and_result125[203]^and_result125[204]^and_result125[205]^and_result125[206]^and_result125[207]^and_result125[208]^and_result125[209]^and_result125[210]^and_result125[211]^and_result125[212]^and_result125[213]^and_result125[214]^and_result125[215]^and_result125[216]^and_result125[217]^and_result125[218]^and_result125[219]^and_result125[220]^and_result125[221]^and_result125[222]^and_result125[223]^and_result125[224]^and_result125[225]^and_result125[226]^and_result125[227]^and_result125[228]^and_result125[229]^and_result125[230]^and_result125[231]^and_result125[232]^and_result125[233]^and_result125[234]^and_result125[235]^and_result125[236]^and_result125[237]^and_result125[238]^and_result125[239]^and_result125[240]^and_result125[241]^and_result125[242]^and_result125[243]^and_result125[244]^and_result125[245]^and_result125[246]^and_result125[247]^and_result125[248]^and_result125[249]^and_result125[250]^and_result125[251]^and_result125[252]^and_result125[253]^and_result125[254];
assign key[126]=and_result126[0]^and_result126[1]^and_result126[2]^and_result126[3]^and_result126[4]^and_result126[5]^and_result126[6]^and_result126[7]^and_result126[8]^and_result126[9]^and_result126[10]^and_result126[11]^and_result126[12]^and_result126[13]^and_result126[14]^and_result126[15]^and_result126[16]^and_result126[17]^and_result126[18]^and_result126[19]^and_result126[20]^and_result126[21]^and_result126[22]^and_result126[23]^and_result126[24]^and_result126[25]^and_result126[26]^and_result126[27]^and_result126[28]^and_result126[29]^and_result126[30]^and_result126[31]^and_result126[32]^and_result126[33]^and_result126[34]^and_result126[35]^and_result126[36]^and_result126[37]^and_result126[38]^and_result126[39]^and_result126[40]^and_result126[41]^and_result126[42]^and_result126[43]^and_result126[44]^and_result126[45]^and_result126[46]^and_result126[47]^and_result126[48]^and_result126[49]^and_result126[50]^and_result126[51]^and_result126[52]^and_result126[53]^and_result126[54]^and_result126[55]^and_result126[56]^and_result126[57]^and_result126[58]^and_result126[59]^and_result126[60]^and_result126[61]^and_result126[62]^and_result126[63]^and_result126[64]^and_result126[65]^and_result126[66]^and_result126[67]^and_result126[68]^and_result126[69]^and_result126[70]^and_result126[71]^and_result126[72]^and_result126[73]^and_result126[74]^and_result126[75]^and_result126[76]^and_result126[77]^and_result126[78]^and_result126[79]^and_result126[80]^and_result126[81]^and_result126[82]^and_result126[83]^and_result126[84]^and_result126[85]^and_result126[86]^and_result126[87]^and_result126[88]^and_result126[89]^and_result126[90]^and_result126[91]^and_result126[92]^and_result126[93]^and_result126[94]^and_result126[95]^and_result126[96]^and_result126[97]^and_result126[98]^and_result126[99]^and_result126[100]^and_result126[101]^and_result126[102]^and_result126[103]^and_result126[104]^and_result126[105]^and_result126[106]^and_result126[107]^and_result126[108]^and_result126[109]^and_result126[110]^and_result126[111]^and_result126[112]^and_result126[113]^and_result126[114]^and_result126[115]^and_result126[116]^and_result126[117]^and_result126[118]^and_result126[119]^and_result126[120]^and_result126[121]^and_result126[122]^and_result126[123]^and_result126[124]^and_result126[125]^and_result126[126]^and_result126[127]^and_result126[128]^and_result126[129]^and_result126[130]^and_result126[131]^and_result126[132]^and_result126[133]^and_result126[134]^and_result126[135]^and_result126[136]^and_result126[137]^and_result126[138]^and_result126[139]^and_result126[140]^and_result126[141]^and_result126[142]^and_result126[143]^and_result126[144]^and_result126[145]^and_result126[146]^and_result126[147]^and_result126[148]^and_result126[149]^and_result126[150]^and_result126[151]^and_result126[152]^and_result126[153]^and_result126[154]^and_result126[155]^and_result126[156]^and_result126[157]^and_result126[158]^and_result126[159]^and_result126[160]^and_result126[161]^and_result126[162]^and_result126[163]^and_result126[164]^and_result126[165]^and_result126[166]^and_result126[167]^and_result126[168]^and_result126[169]^and_result126[170]^and_result126[171]^and_result126[172]^and_result126[173]^and_result126[174]^and_result126[175]^and_result126[176]^and_result126[177]^and_result126[178]^and_result126[179]^and_result126[180]^and_result126[181]^and_result126[182]^and_result126[183]^and_result126[184]^and_result126[185]^and_result126[186]^and_result126[187]^and_result126[188]^and_result126[189]^and_result126[190]^and_result126[191]^and_result126[192]^and_result126[193]^and_result126[194]^and_result126[195]^and_result126[196]^and_result126[197]^and_result126[198]^and_result126[199]^and_result126[200]^and_result126[201]^and_result126[202]^and_result126[203]^and_result126[204]^and_result126[205]^and_result126[206]^and_result126[207]^and_result126[208]^and_result126[209]^and_result126[210]^and_result126[211]^and_result126[212]^and_result126[213]^and_result126[214]^and_result126[215]^and_result126[216]^and_result126[217]^and_result126[218]^and_result126[219]^and_result126[220]^and_result126[221]^and_result126[222]^and_result126[223]^and_result126[224]^and_result126[225]^and_result126[226]^and_result126[227]^and_result126[228]^and_result126[229]^and_result126[230]^and_result126[231]^and_result126[232]^and_result126[233]^and_result126[234]^and_result126[235]^and_result126[236]^and_result126[237]^and_result126[238]^and_result126[239]^and_result126[240]^and_result126[241]^and_result126[242]^and_result126[243]^and_result126[244]^and_result126[245]^and_result126[246]^and_result126[247]^and_result126[248]^and_result126[249]^and_result126[250]^and_result126[251]^and_result126[252]^and_result126[253]^and_result126[254];
assign key[127]=and_result127[0]^and_result127[1]^and_result127[2]^and_result127[3]^and_result127[4]^and_result127[5]^and_result127[6]^and_result127[7]^and_result127[8]^and_result127[9]^and_result127[10]^and_result127[11]^and_result127[12]^and_result127[13]^and_result127[14]^and_result127[15]^and_result127[16]^and_result127[17]^and_result127[18]^and_result127[19]^and_result127[20]^and_result127[21]^and_result127[22]^and_result127[23]^and_result127[24]^and_result127[25]^and_result127[26]^and_result127[27]^and_result127[28]^and_result127[29]^and_result127[30]^and_result127[31]^and_result127[32]^and_result127[33]^and_result127[34]^and_result127[35]^and_result127[36]^and_result127[37]^and_result127[38]^and_result127[39]^and_result127[40]^and_result127[41]^and_result127[42]^and_result127[43]^and_result127[44]^and_result127[45]^and_result127[46]^and_result127[47]^and_result127[48]^and_result127[49]^and_result127[50]^and_result127[51]^and_result127[52]^and_result127[53]^and_result127[54]^and_result127[55]^and_result127[56]^and_result127[57]^and_result127[58]^and_result127[59]^and_result127[60]^and_result127[61]^and_result127[62]^and_result127[63]^and_result127[64]^and_result127[65]^and_result127[66]^and_result127[67]^and_result127[68]^and_result127[69]^and_result127[70]^and_result127[71]^and_result127[72]^and_result127[73]^and_result127[74]^and_result127[75]^and_result127[76]^and_result127[77]^and_result127[78]^and_result127[79]^and_result127[80]^and_result127[81]^and_result127[82]^and_result127[83]^and_result127[84]^and_result127[85]^and_result127[86]^and_result127[87]^and_result127[88]^and_result127[89]^and_result127[90]^and_result127[91]^and_result127[92]^and_result127[93]^and_result127[94]^and_result127[95]^and_result127[96]^and_result127[97]^and_result127[98]^and_result127[99]^and_result127[100]^and_result127[101]^and_result127[102]^and_result127[103]^and_result127[104]^and_result127[105]^and_result127[106]^and_result127[107]^and_result127[108]^and_result127[109]^and_result127[110]^and_result127[111]^and_result127[112]^and_result127[113]^and_result127[114]^and_result127[115]^and_result127[116]^and_result127[117]^and_result127[118]^and_result127[119]^and_result127[120]^and_result127[121]^and_result127[122]^and_result127[123]^and_result127[124]^and_result127[125]^and_result127[126]^and_result127[127]^and_result127[128]^and_result127[129]^and_result127[130]^and_result127[131]^and_result127[132]^and_result127[133]^and_result127[134]^and_result127[135]^and_result127[136]^and_result127[137]^and_result127[138]^and_result127[139]^and_result127[140]^and_result127[141]^and_result127[142]^and_result127[143]^and_result127[144]^and_result127[145]^and_result127[146]^and_result127[147]^and_result127[148]^and_result127[149]^and_result127[150]^and_result127[151]^and_result127[152]^and_result127[153]^and_result127[154]^and_result127[155]^and_result127[156]^and_result127[157]^and_result127[158]^and_result127[159]^and_result127[160]^and_result127[161]^and_result127[162]^and_result127[163]^and_result127[164]^and_result127[165]^and_result127[166]^and_result127[167]^and_result127[168]^and_result127[169]^and_result127[170]^and_result127[171]^and_result127[172]^and_result127[173]^and_result127[174]^and_result127[175]^and_result127[176]^and_result127[177]^and_result127[178]^and_result127[179]^and_result127[180]^and_result127[181]^and_result127[182]^and_result127[183]^and_result127[184]^and_result127[185]^and_result127[186]^and_result127[187]^and_result127[188]^and_result127[189]^and_result127[190]^and_result127[191]^and_result127[192]^and_result127[193]^and_result127[194]^and_result127[195]^and_result127[196]^and_result127[197]^and_result127[198]^and_result127[199]^and_result127[200]^and_result127[201]^and_result127[202]^and_result127[203]^and_result127[204]^and_result127[205]^and_result127[206]^and_result127[207]^and_result127[208]^and_result127[209]^and_result127[210]^and_result127[211]^and_result127[212]^and_result127[213]^and_result127[214]^and_result127[215]^and_result127[216]^and_result127[217]^and_result127[218]^and_result127[219]^and_result127[220]^and_result127[221]^and_result127[222]^and_result127[223]^and_result127[224]^and_result127[225]^and_result127[226]^and_result127[227]^and_result127[228]^and_result127[229]^and_result127[230]^and_result127[231]^and_result127[232]^and_result127[233]^and_result127[234]^and_result127[235]^and_result127[236]^and_result127[237]^and_result127[238]^and_result127[239]^and_result127[240]^and_result127[241]^and_result127[242]^and_result127[243]^and_result127[244]^and_result127[245]^and_result127[246]^and_result127[247]^and_result127[248]^and_result127[249]^and_result127[250]^and_result127[251]^and_result127[252]^and_result127[253]^and_result127[254];
assign key[128]=and_result128[0]^and_result128[1]^and_result128[2]^and_result128[3]^and_result128[4]^and_result128[5]^and_result128[6]^and_result128[7]^and_result128[8]^and_result128[9]^and_result128[10]^and_result128[11]^and_result128[12]^and_result128[13]^and_result128[14]^and_result128[15]^and_result128[16]^and_result128[17]^and_result128[18]^and_result128[19]^and_result128[20]^and_result128[21]^and_result128[22]^and_result128[23]^and_result128[24]^and_result128[25]^and_result128[26]^and_result128[27]^and_result128[28]^and_result128[29]^and_result128[30]^and_result128[31]^and_result128[32]^and_result128[33]^and_result128[34]^and_result128[35]^and_result128[36]^and_result128[37]^and_result128[38]^and_result128[39]^and_result128[40]^and_result128[41]^and_result128[42]^and_result128[43]^and_result128[44]^and_result128[45]^and_result128[46]^and_result128[47]^and_result128[48]^and_result128[49]^and_result128[50]^and_result128[51]^and_result128[52]^and_result128[53]^and_result128[54]^and_result128[55]^and_result128[56]^and_result128[57]^and_result128[58]^and_result128[59]^and_result128[60]^and_result128[61]^and_result128[62]^and_result128[63]^and_result128[64]^and_result128[65]^and_result128[66]^and_result128[67]^and_result128[68]^and_result128[69]^and_result128[70]^and_result128[71]^and_result128[72]^and_result128[73]^and_result128[74]^and_result128[75]^and_result128[76]^and_result128[77]^and_result128[78]^and_result128[79]^and_result128[80]^and_result128[81]^and_result128[82]^and_result128[83]^and_result128[84]^and_result128[85]^and_result128[86]^and_result128[87]^and_result128[88]^and_result128[89]^and_result128[90]^and_result128[91]^and_result128[92]^and_result128[93]^and_result128[94]^and_result128[95]^and_result128[96]^and_result128[97]^and_result128[98]^and_result128[99]^and_result128[100]^and_result128[101]^and_result128[102]^and_result128[103]^and_result128[104]^and_result128[105]^and_result128[106]^and_result128[107]^and_result128[108]^and_result128[109]^and_result128[110]^and_result128[111]^and_result128[112]^and_result128[113]^and_result128[114]^and_result128[115]^and_result128[116]^and_result128[117]^and_result128[118]^and_result128[119]^and_result128[120]^and_result128[121]^and_result128[122]^and_result128[123]^and_result128[124]^and_result128[125]^and_result128[126]^and_result128[127]^and_result128[128]^and_result128[129]^and_result128[130]^and_result128[131]^and_result128[132]^and_result128[133]^and_result128[134]^and_result128[135]^and_result128[136]^and_result128[137]^and_result128[138]^and_result128[139]^and_result128[140]^and_result128[141]^and_result128[142]^and_result128[143]^and_result128[144]^and_result128[145]^and_result128[146]^and_result128[147]^and_result128[148]^and_result128[149]^and_result128[150]^and_result128[151]^and_result128[152]^and_result128[153]^and_result128[154]^and_result128[155]^and_result128[156]^and_result128[157]^and_result128[158]^and_result128[159]^and_result128[160]^and_result128[161]^and_result128[162]^and_result128[163]^and_result128[164]^and_result128[165]^and_result128[166]^and_result128[167]^and_result128[168]^and_result128[169]^and_result128[170]^and_result128[171]^and_result128[172]^and_result128[173]^and_result128[174]^and_result128[175]^and_result128[176]^and_result128[177]^and_result128[178]^and_result128[179]^and_result128[180]^and_result128[181]^and_result128[182]^and_result128[183]^and_result128[184]^and_result128[185]^and_result128[186]^and_result128[187]^and_result128[188]^and_result128[189]^and_result128[190]^and_result128[191]^and_result128[192]^and_result128[193]^and_result128[194]^and_result128[195]^and_result128[196]^and_result128[197]^and_result128[198]^and_result128[199]^and_result128[200]^and_result128[201]^and_result128[202]^and_result128[203]^and_result128[204]^and_result128[205]^and_result128[206]^and_result128[207]^and_result128[208]^and_result128[209]^and_result128[210]^and_result128[211]^and_result128[212]^and_result128[213]^and_result128[214]^and_result128[215]^and_result128[216]^and_result128[217]^and_result128[218]^and_result128[219]^and_result128[220]^and_result128[221]^and_result128[222]^and_result128[223]^and_result128[224]^and_result128[225]^and_result128[226]^and_result128[227]^and_result128[228]^and_result128[229]^and_result128[230]^and_result128[231]^and_result128[232]^and_result128[233]^and_result128[234]^and_result128[235]^and_result128[236]^and_result128[237]^and_result128[238]^and_result128[239]^and_result128[240]^and_result128[241]^and_result128[242]^and_result128[243]^and_result128[244]^and_result128[245]^and_result128[246]^and_result128[247]^and_result128[248]^and_result128[249]^and_result128[250]^and_result128[251]^and_result128[252]^and_result128[253]^and_result128[254];
assign key[129]=and_result129[0]^and_result129[1]^and_result129[2]^and_result129[3]^and_result129[4]^and_result129[5]^and_result129[6]^and_result129[7]^and_result129[8]^and_result129[9]^and_result129[10]^and_result129[11]^and_result129[12]^and_result129[13]^and_result129[14]^and_result129[15]^and_result129[16]^and_result129[17]^and_result129[18]^and_result129[19]^and_result129[20]^and_result129[21]^and_result129[22]^and_result129[23]^and_result129[24]^and_result129[25]^and_result129[26]^and_result129[27]^and_result129[28]^and_result129[29]^and_result129[30]^and_result129[31]^and_result129[32]^and_result129[33]^and_result129[34]^and_result129[35]^and_result129[36]^and_result129[37]^and_result129[38]^and_result129[39]^and_result129[40]^and_result129[41]^and_result129[42]^and_result129[43]^and_result129[44]^and_result129[45]^and_result129[46]^and_result129[47]^and_result129[48]^and_result129[49]^and_result129[50]^and_result129[51]^and_result129[52]^and_result129[53]^and_result129[54]^and_result129[55]^and_result129[56]^and_result129[57]^and_result129[58]^and_result129[59]^and_result129[60]^and_result129[61]^and_result129[62]^and_result129[63]^and_result129[64]^and_result129[65]^and_result129[66]^and_result129[67]^and_result129[68]^and_result129[69]^and_result129[70]^and_result129[71]^and_result129[72]^and_result129[73]^and_result129[74]^and_result129[75]^and_result129[76]^and_result129[77]^and_result129[78]^and_result129[79]^and_result129[80]^and_result129[81]^and_result129[82]^and_result129[83]^and_result129[84]^and_result129[85]^and_result129[86]^and_result129[87]^and_result129[88]^and_result129[89]^and_result129[90]^and_result129[91]^and_result129[92]^and_result129[93]^and_result129[94]^and_result129[95]^and_result129[96]^and_result129[97]^and_result129[98]^and_result129[99]^and_result129[100]^and_result129[101]^and_result129[102]^and_result129[103]^and_result129[104]^and_result129[105]^and_result129[106]^and_result129[107]^and_result129[108]^and_result129[109]^and_result129[110]^and_result129[111]^and_result129[112]^and_result129[113]^and_result129[114]^and_result129[115]^and_result129[116]^and_result129[117]^and_result129[118]^and_result129[119]^and_result129[120]^and_result129[121]^and_result129[122]^and_result129[123]^and_result129[124]^and_result129[125]^and_result129[126]^and_result129[127]^and_result129[128]^and_result129[129]^and_result129[130]^and_result129[131]^and_result129[132]^and_result129[133]^and_result129[134]^and_result129[135]^and_result129[136]^and_result129[137]^and_result129[138]^and_result129[139]^and_result129[140]^and_result129[141]^and_result129[142]^and_result129[143]^and_result129[144]^and_result129[145]^and_result129[146]^and_result129[147]^and_result129[148]^and_result129[149]^and_result129[150]^and_result129[151]^and_result129[152]^and_result129[153]^and_result129[154]^and_result129[155]^and_result129[156]^and_result129[157]^and_result129[158]^and_result129[159]^and_result129[160]^and_result129[161]^and_result129[162]^and_result129[163]^and_result129[164]^and_result129[165]^and_result129[166]^and_result129[167]^and_result129[168]^and_result129[169]^and_result129[170]^and_result129[171]^and_result129[172]^and_result129[173]^and_result129[174]^and_result129[175]^and_result129[176]^and_result129[177]^and_result129[178]^and_result129[179]^and_result129[180]^and_result129[181]^and_result129[182]^and_result129[183]^and_result129[184]^and_result129[185]^and_result129[186]^and_result129[187]^and_result129[188]^and_result129[189]^and_result129[190]^and_result129[191]^and_result129[192]^and_result129[193]^and_result129[194]^and_result129[195]^and_result129[196]^and_result129[197]^and_result129[198]^and_result129[199]^and_result129[200]^and_result129[201]^and_result129[202]^and_result129[203]^and_result129[204]^and_result129[205]^and_result129[206]^and_result129[207]^and_result129[208]^and_result129[209]^and_result129[210]^and_result129[211]^and_result129[212]^and_result129[213]^and_result129[214]^and_result129[215]^and_result129[216]^and_result129[217]^and_result129[218]^and_result129[219]^and_result129[220]^and_result129[221]^and_result129[222]^and_result129[223]^and_result129[224]^and_result129[225]^and_result129[226]^and_result129[227]^and_result129[228]^and_result129[229]^and_result129[230]^and_result129[231]^and_result129[232]^and_result129[233]^and_result129[234]^and_result129[235]^and_result129[236]^and_result129[237]^and_result129[238]^and_result129[239]^and_result129[240]^and_result129[241]^and_result129[242]^and_result129[243]^and_result129[244]^and_result129[245]^and_result129[246]^and_result129[247]^and_result129[248]^and_result129[249]^and_result129[250]^and_result129[251]^and_result129[252]^and_result129[253]^and_result129[254];
assign key[130]=and_result130[0]^and_result130[1]^and_result130[2]^and_result130[3]^and_result130[4]^and_result130[5]^and_result130[6]^and_result130[7]^and_result130[8]^and_result130[9]^and_result130[10]^and_result130[11]^and_result130[12]^and_result130[13]^and_result130[14]^and_result130[15]^and_result130[16]^and_result130[17]^and_result130[18]^and_result130[19]^and_result130[20]^and_result130[21]^and_result130[22]^and_result130[23]^and_result130[24]^and_result130[25]^and_result130[26]^and_result130[27]^and_result130[28]^and_result130[29]^and_result130[30]^and_result130[31]^and_result130[32]^and_result130[33]^and_result130[34]^and_result130[35]^and_result130[36]^and_result130[37]^and_result130[38]^and_result130[39]^and_result130[40]^and_result130[41]^and_result130[42]^and_result130[43]^and_result130[44]^and_result130[45]^and_result130[46]^and_result130[47]^and_result130[48]^and_result130[49]^and_result130[50]^and_result130[51]^and_result130[52]^and_result130[53]^and_result130[54]^and_result130[55]^and_result130[56]^and_result130[57]^and_result130[58]^and_result130[59]^and_result130[60]^and_result130[61]^and_result130[62]^and_result130[63]^and_result130[64]^and_result130[65]^and_result130[66]^and_result130[67]^and_result130[68]^and_result130[69]^and_result130[70]^and_result130[71]^and_result130[72]^and_result130[73]^and_result130[74]^and_result130[75]^and_result130[76]^and_result130[77]^and_result130[78]^and_result130[79]^and_result130[80]^and_result130[81]^and_result130[82]^and_result130[83]^and_result130[84]^and_result130[85]^and_result130[86]^and_result130[87]^and_result130[88]^and_result130[89]^and_result130[90]^and_result130[91]^and_result130[92]^and_result130[93]^and_result130[94]^and_result130[95]^and_result130[96]^and_result130[97]^and_result130[98]^and_result130[99]^and_result130[100]^and_result130[101]^and_result130[102]^and_result130[103]^and_result130[104]^and_result130[105]^and_result130[106]^and_result130[107]^and_result130[108]^and_result130[109]^and_result130[110]^and_result130[111]^and_result130[112]^and_result130[113]^and_result130[114]^and_result130[115]^and_result130[116]^and_result130[117]^and_result130[118]^and_result130[119]^and_result130[120]^and_result130[121]^and_result130[122]^and_result130[123]^and_result130[124]^and_result130[125]^and_result130[126]^and_result130[127]^and_result130[128]^and_result130[129]^and_result130[130]^and_result130[131]^and_result130[132]^and_result130[133]^and_result130[134]^and_result130[135]^and_result130[136]^and_result130[137]^and_result130[138]^and_result130[139]^and_result130[140]^and_result130[141]^and_result130[142]^and_result130[143]^and_result130[144]^and_result130[145]^and_result130[146]^and_result130[147]^and_result130[148]^and_result130[149]^and_result130[150]^and_result130[151]^and_result130[152]^and_result130[153]^and_result130[154]^and_result130[155]^and_result130[156]^and_result130[157]^and_result130[158]^and_result130[159]^and_result130[160]^and_result130[161]^and_result130[162]^and_result130[163]^and_result130[164]^and_result130[165]^and_result130[166]^and_result130[167]^and_result130[168]^and_result130[169]^and_result130[170]^and_result130[171]^and_result130[172]^and_result130[173]^and_result130[174]^and_result130[175]^and_result130[176]^and_result130[177]^and_result130[178]^and_result130[179]^and_result130[180]^and_result130[181]^and_result130[182]^and_result130[183]^and_result130[184]^and_result130[185]^and_result130[186]^and_result130[187]^and_result130[188]^and_result130[189]^and_result130[190]^and_result130[191]^and_result130[192]^and_result130[193]^and_result130[194]^and_result130[195]^and_result130[196]^and_result130[197]^and_result130[198]^and_result130[199]^and_result130[200]^and_result130[201]^and_result130[202]^and_result130[203]^and_result130[204]^and_result130[205]^and_result130[206]^and_result130[207]^and_result130[208]^and_result130[209]^and_result130[210]^and_result130[211]^and_result130[212]^and_result130[213]^and_result130[214]^and_result130[215]^and_result130[216]^and_result130[217]^and_result130[218]^and_result130[219]^and_result130[220]^and_result130[221]^and_result130[222]^and_result130[223]^and_result130[224]^and_result130[225]^and_result130[226]^and_result130[227]^and_result130[228]^and_result130[229]^and_result130[230]^and_result130[231]^and_result130[232]^and_result130[233]^and_result130[234]^and_result130[235]^and_result130[236]^and_result130[237]^and_result130[238]^and_result130[239]^and_result130[240]^and_result130[241]^and_result130[242]^and_result130[243]^and_result130[244]^and_result130[245]^and_result130[246]^and_result130[247]^and_result130[248]^and_result130[249]^and_result130[250]^and_result130[251]^and_result130[252]^and_result130[253]^and_result130[254];
assign key[131]=and_result131[0]^and_result131[1]^and_result131[2]^and_result131[3]^and_result131[4]^and_result131[5]^and_result131[6]^and_result131[7]^and_result131[8]^and_result131[9]^and_result131[10]^and_result131[11]^and_result131[12]^and_result131[13]^and_result131[14]^and_result131[15]^and_result131[16]^and_result131[17]^and_result131[18]^and_result131[19]^and_result131[20]^and_result131[21]^and_result131[22]^and_result131[23]^and_result131[24]^and_result131[25]^and_result131[26]^and_result131[27]^and_result131[28]^and_result131[29]^and_result131[30]^and_result131[31]^and_result131[32]^and_result131[33]^and_result131[34]^and_result131[35]^and_result131[36]^and_result131[37]^and_result131[38]^and_result131[39]^and_result131[40]^and_result131[41]^and_result131[42]^and_result131[43]^and_result131[44]^and_result131[45]^and_result131[46]^and_result131[47]^and_result131[48]^and_result131[49]^and_result131[50]^and_result131[51]^and_result131[52]^and_result131[53]^and_result131[54]^and_result131[55]^and_result131[56]^and_result131[57]^and_result131[58]^and_result131[59]^and_result131[60]^and_result131[61]^and_result131[62]^and_result131[63]^and_result131[64]^and_result131[65]^and_result131[66]^and_result131[67]^and_result131[68]^and_result131[69]^and_result131[70]^and_result131[71]^and_result131[72]^and_result131[73]^and_result131[74]^and_result131[75]^and_result131[76]^and_result131[77]^and_result131[78]^and_result131[79]^and_result131[80]^and_result131[81]^and_result131[82]^and_result131[83]^and_result131[84]^and_result131[85]^and_result131[86]^and_result131[87]^and_result131[88]^and_result131[89]^and_result131[90]^and_result131[91]^and_result131[92]^and_result131[93]^and_result131[94]^and_result131[95]^and_result131[96]^and_result131[97]^and_result131[98]^and_result131[99]^and_result131[100]^and_result131[101]^and_result131[102]^and_result131[103]^and_result131[104]^and_result131[105]^and_result131[106]^and_result131[107]^and_result131[108]^and_result131[109]^and_result131[110]^and_result131[111]^and_result131[112]^and_result131[113]^and_result131[114]^and_result131[115]^and_result131[116]^and_result131[117]^and_result131[118]^and_result131[119]^and_result131[120]^and_result131[121]^and_result131[122]^and_result131[123]^and_result131[124]^and_result131[125]^and_result131[126]^and_result131[127]^and_result131[128]^and_result131[129]^and_result131[130]^and_result131[131]^and_result131[132]^and_result131[133]^and_result131[134]^and_result131[135]^and_result131[136]^and_result131[137]^and_result131[138]^and_result131[139]^and_result131[140]^and_result131[141]^and_result131[142]^and_result131[143]^and_result131[144]^and_result131[145]^and_result131[146]^and_result131[147]^and_result131[148]^and_result131[149]^and_result131[150]^and_result131[151]^and_result131[152]^and_result131[153]^and_result131[154]^and_result131[155]^and_result131[156]^and_result131[157]^and_result131[158]^and_result131[159]^and_result131[160]^and_result131[161]^and_result131[162]^and_result131[163]^and_result131[164]^and_result131[165]^and_result131[166]^and_result131[167]^and_result131[168]^and_result131[169]^and_result131[170]^and_result131[171]^and_result131[172]^and_result131[173]^and_result131[174]^and_result131[175]^and_result131[176]^and_result131[177]^and_result131[178]^and_result131[179]^and_result131[180]^and_result131[181]^and_result131[182]^and_result131[183]^and_result131[184]^and_result131[185]^and_result131[186]^and_result131[187]^and_result131[188]^and_result131[189]^and_result131[190]^and_result131[191]^and_result131[192]^and_result131[193]^and_result131[194]^and_result131[195]^and_result131[196]^and_result131[197]^and_result131[198]^and_result131[199]^and_result131[200]^and_result131[201]^and_result131[202]^and_result131[203]^and_result131[204]^and_result131[205]^and_result131[206]^and_result131[207]^and_result131[208]^and_result131[209]^and_result131[210]^and_result131[211]^and_result131[212]^and_result131[213]^and_result131[214]^and_result131[215]^and_result131[216]^and_result131[217]^and_result131[218]^and_result131[219]^and_result131[220]^and_result131[221]^and_result131[222]^and_result131[223]^and_result131[224]^and_result131[225]^and_result131[226]^and_result131[227]^and_result131[228]^and_result131[229]^and_result131[230]^and_result131[231]^and_result131[232]^and_result131[233]^and_result131[234]^and_result131[235]^and_result131[236]^and_result131[237]^and_result131[238]^and_result131[239]^and_result131[240]^and_result131[241]^and_result131[242]^and_result131[243]^and_result131[244]^and_result131[245]^and_result131[246]^and_result131[247]^and_result131[248]^and_result131[249]^and_result131[250]^and_result131[251]^and_result131[252]^and_result131[253]^and_result131[254];
assign key[132]=and_result132[0]^and_result132[1]^and_result132[2]^and_result132[3]^and_result132[4]^and_result132[5]^and_result132[6]^and_result132[7]^and_result132[8]^and_result132[9]^and_result132[10]^and_result132[11]^and_result132[12]^and_result132[13]^and_result132[14]^and_result132[15]^and_result132[16]^and_result132[17]^and_result132[18]^and_result132[19]^and_result132[20]^and_result132[21]^and_result132[22]^and_result132[23]^and_result132[24]^and_result132[25]^and_result132[26]^and_result132[27]^and_result132[28]^and_result132[29]^and_result132[30]^and_result132[31]^and_result132[32]^and_result132[33]^and_result132[34]^and_result132[35]^and_result132[36]^and_result132[37]^and_result132[38]^and_result132[39]^and_result132[40]^and_result132[41]^and_result132[42]^and_result132[43]^and_result132[44]^and_result132[45]^and_result132[46]^and_result132[47]^and_result132[48]^and_result132[49]^and_result132[50]^and_result132[51]^and_result132[52]^and_result132[53]^and_result132[54]^and_result132[55]^and_result132[56]^and_result132[57]^and_result132[58]^and_result132[59]^and_result132[60]^and_result132[61]^and_result132[62]^and_result132[63]^and_result132[64]^and_result132[65]^and_result132[66]^and_result132[67]^and_result132[68]^and_result132[69]^and_result132[70]^and_result132[71]^and_result132[72]^and_result132[73]^and_result132[74]^and_result132[75]^and_result132[76]^and_result132[77]^and_result132[78]^and_result132[79]^and_result132[80]^and_result132[81]^and_result132[82]^and_result132[83]^and_result132[84]^and_result132[85]^and_result132[86]^and_result132[87]^and_result132[88]^and_result132[89]^and_result132[90]^and_result132[91]^and_result132[92]^and_result132[93]^and_result132[94]^and_result132[95]^and_result132[96]^and_result132[97]^and_result132[98]^and_result132[99]^and_result132[100]^and_result132[101]^and_result132[102]^and_result132[103]^and_result132[104]^and_result132[105]^and_result132[106]^and_result132[107]^and_result132[108]^and_result132[109]^and_result132[110]^and_result132[111]^and_result132[112]^and_result132[113]^and_result132[114]^and_result132[115]^and_result132[116]^and_result132[117]^and_result132[118]^and_result132[119]^and_result132[120]^and_result132[121]^and_result132[122]^and_result132[123]^and_result132[124]^and_result132[125]^and_result132[126]^and_result132[127]^and_result132[128]^and_result132[129]^and_result132[130]^and_result132[131]^and_result132[132]^and_result132[133]^and_result132[134]^and_result132[135]^and_result132[136]^and_result132[137]^and_result132[138]^and_result132[139]^and_result132[140]^and_result132[141]^and_result132[142]^and_result132[143]^and_result132[144]^and_result132[145]^and_result132[146]^and_result132[147]^and_result132[148]^and_result132[149]^and_result132[150]^and_result132[151]^and_result132[152]^and_result132[153]^and_result132[154]^and_result132[155]^and_result132[156]^and_result132[157]^and_result132[158]^and_result132[159]^and_result132[160]^and_result132[161]^and_result132[162]^and_result132[163]^and_result132[164]^and_result132[165]^and_result132[166]^and_result132[167]^and_result132[168]^and_result132[169]^and_result132[170]^and_result132[171]^and_result132[172]^and_result132[173]^and_result132[174]^and_result132[175]^and_result132[176]^and_result132[177]^and_result132[178]^and_result132[179]^and_result132[180]^and_result132[181]^and_result132[182]^and_result132[183]^and_result132[184]^and_result132[185]^and_result132[186]^and_result132[187]^and_result132[188]^and_result132[189]^and_result132[190]^and_result132[191]^and_result132[192]^and_result132[193]^and_result132[194]^and_result132[195]^and_result132[196]^and_result132[197]^and_result132[198]^and_result132[199]^and_result132[200]^and_result132[201]^and_result132[202]^and_result132[203]^and_result132[204]^and_result132[205]^and_result132[206]^and_result132[207]^and_result132[208]^and_result132[209]^and_result132[210]^and_result132[211]^and_result132[212]^and_result132[213]^and_result132[214]^and_result132[215]^and_result132[216]^and_result132[217]^and_result132[218]^and_result132[219]^and_result132[220]^and_result132[221]^and_result132[222]^and_result132[223]^and_result132[224]^and_result132[225]^and_result132[226]^and_result132[227]^and_result132[228]^and_result132[229]^and_result132[230]^and_result132[231]^and_result132[232]^and_result132[233]^and_result132[234]^and_result132[235]^and_result132[236]^and_result132[237]^and_result132[238]^and_result132[239]^and_result132[240]^and_result132[241]^and_result132[242]^and_result132[243]^and_result132[244]^and_result132[245]^and_result132[246]^and_result132[247]^and_result132[248]^and_result132[249]^and_result132[250]^and_result132[251]^and_result132[252]^and_result132[253]^and_result132[254];
assign key[133]=and_result133[0]^and_result133[1]^and_result133[2]^and_result133[3]^and_result133[4]^and_result133[5]^and_result133[6]^and_result133[7]^and_result133[8]^and_result133[9]^and_result133[10]^and_result133[11]^and_result133[12]^and_result133[13]^and_result133[14]^and_result133[15]^and_result133[16]^and_result133[17]^and_result133[18]^and_result133[19]^and_result133[20]^and_result133[21]^and_result133[22]^and_result133[23]^and_result133[24]^and_result133[25]^and_result133[26]^and_result133[27]^and_result133[28]^and_result133[29]^and_result133[30]^and_result133[31]^and_result133[32]^and_result133[33]^and_result133[34]^and_result133[35]^and_result133[36]^and_result133[37]^and_result133[38]^and_result133[39]^and_result133[40]^and_result133[41]^and_result133[42]^and_result133[43]^and_result133[44]^and_result133[45]^and_result133[46]^and_result133[47]^and_result133[48]^and_result133[49]^and_result133[50]^and_result133[51]^and_result133[52]^and_result133[53]^and_result133[54]^and_result133[55]^and_result133[56]^and_result133[57]^and_result133[58]^and_result133[59]^and_result133[60]^and_result133[61]^and_result133[62]^and_result133[63]^and_result133[64]^and_result133[65]^and_result133[66]^and_result133[67]^and_result133[68]^and_result133[69]^and_result133[70]^and_result133[71]^and_result133[72]^and_result133[73]^and_result133[74]^and_result133[75]^and_result133[76]^and_result133[77]^and_result133[78]^and_result133[79]^and_result133[80]^and_result133[81]^and_result133[82]^and_result133[83]^and_result133[84]^and_result133[85]^and_result133[86]^and_result133[87]^and_result133[88]^and_result133[89]^and_result133[90]^and_result133[91]^and_result133[92]^and_result133[93]^and_result133[94]^and_result133[95]^and_result133[96]^and_result133[97]^and_result133[98]^and_result133[99]^and_result133[100]^and_result133[101]^and_result133[102]^and_result133[103]^and_result133[104]^and_result133[105]^and_result133[106]^and_result133[107]^and_result133[108]^and_result133[109]^and_result133[110]^and_result133[111]^and_result133[112]^and_result133[113]^and_result133[114]^and_result133[115]^and_result133[116]^and_result133[117]^and_result133[118]^and_result133[119]^and_result133[120]^and_result133[121]^and_result133[122]^and_result133[123]^and_result133[124]^and_result133[125]^and_result133[126]^and_result133[127]^and_result133[128]^and_result133[129]^and_result133[130]^and_result133[131]^and_result133[132]^and_result133[133]^and_result133[134]^and_result133[135]^and_result133[136]^and_result133[137]^and_result133[138]^and_result133[139]^and_result133[140]^and_result133[141]^and_result133[142]^and_result133[143]^and_result133[144]^and_result133[145]^and_result133[146]^and_result133[147]^and_result133[148]^and_result133[149]^and_result133[150]^and_result133[151]^and_result133[152]^and_result133[153]^and_result133[154]^and_result133[155]^and_result133[156]^and_result133[157]^and_result133[158]^and_result133[159]^and_result133[160]^and_result133[161]^and_result133[162]^and_result133[163]^and_result133[164]^and_result133[165]^and_result133[166]^and_result133[167]^and_result133[168]^and_result133[169]^and_result133[170]^and_result133[171]^and_result133[172]^and_result133[173]^and_result133[174]^and_result133[175]^and_result133[176]^and_result133[177]^and_result133[178]^and_result133[179]^and_result133[180]^and_result133[181]^and_result133[182]^and_result133[183]^and_result133[184]^and_result133[185]^and_result133[186]^and_result133[187]^and_result133[188]^and_result133[189]^and_result133[190]^and_result133[191]^and_result133[192]^and_result133[193]^and_result133[194]^and_result133[195]^and_result133[196]^and_result133[197]^and_result133[198]^and_result133[199]^and_result133[200]^and_result133[201]^and_result133[202]^and_result133[203]^and_result133[204]^and_result133[205]^and_result133[206]^and_result133[207]^and_result133[208]^and_result133[209]^and_result133[210]^and_result133[211]^and_result133[212]^and_result133[213]^and_result133[214]^and_result133[215]^and_result133[216]^and_result133[217]^and_result133[218]^and_result133[219]^and_result133[220]^and_result133[221]^and_result133[222]^and_result133[223]^and_result133[224]^and_result133[225]^and_result133[226]^and_result133[227]^and_result133[228]^and_result133[229]^and_result133[230]^and_result133[231]^and_result133[232]^and_result133[233]^and_result133[234]^and_result133[235]^and_result133[236]^and_result133[237]^and_result133[238]^and_result133[239]^and_result133[240]^and_result133[241]^and_result133[242]^and_result133[243]^and_result133[244]^and_result133[245]^and_result133[246]^and_result133[247]^and_result133[248]^and_result133[249]^and_result133[250]^and_result133[251]^and_result133[252]^and_result133[253]^and_result133[254];
assign key[134]=and_result134[0]^and_result134[1]^and_result134[2]^and_result134[3]^and_result134[4]^and_result134[5]^and_result134[6]^and_result134[7]^and_result134[8]^and_result134[9]^and_result134[10]^and_result134[11]^and_result134[12]^and_result134[13]^and_result134[14]^and_result134[15]^and_result134[16]^and_result134[17]^and_result134[18]^and_result134[19]^and_result134[20]^and_result134[21]^and_result134[22]^and_result134[23]^and_result134[24]^and_result134[25]^and_result134[26]^and_result134[27]^and_result134[28]^and_result134[29]^and_result134[30]^and_result134[31]^and_result134[32]^and_result134[33]^and_result134[34]^and_result134[35]^and_result134[36]^and_result134[37]^and_result134[38]^and_result134[39]^and_result134[40]^and_result134[41]^and_result134[42]^and_result134[43]^and_result134[44]^and_result134[45]^and_result134[46]^and_result134[47]^and_result134[48]^and_result134[49]^and_result134[50]^and_result134[51]^and_result134[52]^and_result134[53]^and_result134[54]^and_result134[55]^and_result134[56]^and_result134[57]^and_result134[58]^and_result134[59]^and_result134[60]^and_result134[61]^and_result134[62]^and_result134[63]^and_result134[64]^and_result134[65]^and_result134[66]^and_result134[67]^and_result134[68]^and_result134[69]^and_result134[70]^and_result134[71]^and_result134[72]^and_result134[73]^and_result134[74]^and_result134[75]^and_result134[76]^and_result134[77]^and_result134[78]^and_result134[79]^and_result134[80]^and_result134[81]^and_result134[82]^and_result134[83]^and_result134[84]^and_result134[85]^and_result134[86]^and_result134[87]^and_result134[88]^and_result134[89]^and_result134[90]^and_result134[91]^and_result134[92]^and_result134[93]^and_result134[94]^and_result134[95]^and_result134[96]^and_result134[97]^and_result134[98]^and_result134[99]^and_result134[100]^and_result134[101]^and_result134[102]^and_result134[103]^and_result134[104]^and_result134[105]^and_result134[106]^and_result134[107]^and_result134[108]^and_result134[109]^and_result134[110]^and_result134[111]^and_result134[112]^and_result134[113]^and_result134[114]^and_result134[115]^and_result134[116]^and_result134[117]^and_result134[118]^and_result134[119]^and_result134[120]^and_result134[121]^and_result134[122]^and_result134[123]^and_result134[124]^and_result134[125]^and_result134[126]^and_result134[127]^and_result134[128]^and_result134[129]^and_result134[130]^and_result134[131]^and_result134[132]^and_result134[133]^and_result134[134]^and_result134[135]^and_result134[136]^and_result134[137]^and_result134[138]^and_result134[139]^and_result134[140]^and_result134[141]^and_result134[142]^and_result134[143]^and_result134[144]^and_result134[145]^and_result134[146]^and_result134[147]^and_result134[148]^and_result134[149]^and_result134[150]^and_result134[151]^and_result134[152]^and_result134[153]^and_result134[154]^and_result134[155]^and_result134[156]^and_result134[157]^and_result134[158]^and_result134[159]^and_result134[160]^and_result134[161]^and_result134[162]^and_result134[163]^and_result134[164]^and_result134[165]^and_result134[166]^and_result134[167]^and_result134[168]^and_result134[169]^and_result134[170]^and_result134[171]^and_result134[172]^and_result134[173]^and_result134[174]^and_result134[175]^and_result134[176]^and_result134[177]^and_result134[178]^and_result134[179]^and_result134[180]^and_result134[181]^and_result134[182]^and_result134[183]^and_result134[184]^and_result134[185]^and_result134[186]^and_result134[187]^and_result134[188]^and_result134[189]^and_result134[190]^and_result134[191]^and_result134[192]^and_result134[193]^and_result134[194]^and_result134[195]^and_result134[196]^and_result134[197]^and_result134[198]^and_result134[199]^and_result134[200]^and_result134[201]^and_result134[202]^and_result134[203]^and_result134[204]^and_result134[205]^and_result134[206]^and_result134[207]^and_result134[208]^and_result134[209]^and_result134[210]^and_result134[211]^and_result134[212]^and_result134[213]^and_result134[214]^and_result134[215]^and_result134[216]^and_result134[217]^and_result134[218]^and_result134[219]^and_result134[220]^and_result134[221]^and_result134[222]^and_result134[223]^and_result134[224]^and_result134[225]^and_result134[226]^and_result134[227]^and_result134[228]^and_result134[229]^and_result134[230]^and_result134[231]^and_result134[232]^and_result134[233]^and_result134[234]^and_result134[235]^and_result134[236]^and_result134[237]^and_result134[238]^and_result134[239]^and_result134[240]^and_result134[241]^and_result134[242]^and_result134[243]^and_result134[244]^and_result134[245]^and_result134[246]^and_result134[247]^and_result134[248]^and_result134[249]^and_result134[250]^and_result134[251]^and_result134[252]^and_result134[253]^and_result134[254];
assign key[135]=and_result135[0]^and_result135[1]^and_result135[2]^and_result135[3]^and_result135[4]^and_result135[5]^and_result135[6]^and_result135[7]^and_result135[8]^and_result135[9]^and_result135[10]^and_result135[11]^and_result135[12]^and_result135[13]^and_result135[14]^and_result135[15]^and_result135[16]^and_result135[17]^and_result135[18]^and_result135[19]^and_result135[20]^and_result135[21]^and_result135[22]^and_result135[23]^and_result135[24]^and_result135[25]^and_result135[26]^and_result135[27]^and_result135[28]^and_result135[29]^and_result135[30]^and_result135[31]^and_result135[32]^and_result135[33]^and_result135[34]^and_result135[35]^and_result135[36]^and_result135[37]^and_result135[38]^and_result135[39]^and_result135[40]^and_result135[41]^and_result135[42]^and_result135[43]^and_result135[44]^and_result135[45]^and_result135[46]^and_result135[47]^and_result135[48]^and_result135[49]^and_result135[50]^and_result135[51]^and_result135[52]^and_result135[53]^and_result135[54]^and_result135[55]^and_result135[56]^and_result135[57]^and_result135[58]^and_result135[59]^and_result135[60]^and_result135[61]^and_result135[62]^and_result135[63]^and_result135[64]^and_result135[65]^and_result135[66]^and_result135[67]^and_result135[68]^and_result135[69]^and_result135[70]^and_result135[71]^and_result135[72]^and_result135[73]^and_result135[74]^and_result135[75]^and_result135[76]^and_result135[77]^and_result135[78]^and_result135[79]^and_result135[80]^and_result135[81]^and_result135[82]^and_result135[83]^and_result135[84]^and_result135[85]^and_result135[86]^and_result135[87]^and_result135[88]^and_result135[89]^and_result135[90]^and_result135[91]^and_result135[92]^and_result135[93]^and_result135[94]^and_result135[95]^and_result135[96]^and_result135[97]^and_result135[98]^and_result135[99]^and_result135[100]^and_result135[101]^and_result135[102]^and_result135[103]^and_result135[104]^and_result135[105]^and_result135[106]^and_result135[107]^and_result135[108]^and_result135[109]^and_result135[110]^and_result135[111]^and_result135[112]^and_result135[113]^and_result135[114]^and_result135[115]^and_result135[116]^and_result135[117]^and_result135[118]^and_result135[119]^and_result135[120]^and_result135[121]^and_result135[122]^and_result135[123]^and_result135[124]^and_result135[125]^and_result135[126]^and_result135[127]^and_result135[128]^and_result135[129]^and_result135[130]^and_result135[131]^and_result135[132]^and_result135[133]^and_result135[134]^and_result135[135]^and_result135[136]^and_result135[137]^and_result135[138]^and_result135[139]^and_result135[140]^and_result135[141]^and_result135[142]^and_result135[143]^and_result135[144]^and_result135[145]^and_result135[146]^and_result135[147]^and_result135[148]^and_result135[149]^and_result135[150]^and_result135[151]^and_result135[152]^and_result135[153]^and_result135[154]^and_result135[155]^and_result135[156]^and_result135[157]^and_result135[158]^and_result135[159]^and_result135[160]^and_result135[161]^and_result135[162]^and_result135[163]^and_result135[164]^and_result135[165]^and_result135[166]^and_result135[167]^and_result135[168]^and_result135[169]^and_result135[170]^and_result135[171]^and_result135[172]^and_result135[173]^and_result135[174]^and_result135[175]^and_result135[176]^and_result135[177]^and_result135[178]^and_result135[179]^and_result135[180]^and_result135[181]^and_result135[182]^and_result135[183]^and_result135[184]^and_result135[185]^and_result135[186]^and_result135[187]^and_result135[188]^and_result135[189]^and_result135[190]^and_result135[191]^and_result135[192]^and_result135[193]^and_result135[194]^and_result135[195]^and_result135[196]^and_result135[197]^and_result135[198]^and_result135[199]^and_result135[200]^and_result135[201]^and_result135[202]^and_result135[203]^and_result135[204]^and_result135[205]^and_result135[206]^and_result135[207]^and_result135[208]^and_result135[209]^and_result135[210]^and_result135[211]^and_result135[212]^and_result135[213]^and_result135[214]^and_result135[215]^and_result135[216]^and_result135[217]^and_result135[218]^and_result135[219]^and_result135[220]^and_result135[221]^and_result135[222]^and_result135[223]^and_result135[224]^and_result135[225]^and_result135[226]^and_result135[227]^and_result135[228]^and_result135[229]^and_result135[230]^and_result135[231]^and_result135[232]^and_result135[233]^and_result135[234]^and_result135[235]^and_result135[236]^and_result135[237]^and_result135[238]^and_result135[239]^and_result135[240]^and_result135[241]^and_result135[242]^and_result135[243]^and_result135[244]^and_result135[245]^and_result135[246]^and_result135[247]^and_result135[248]^and_result135[249]^and_result135[250]^and_result135[251]^and_result135[252]^and_result135[253]^and_result135[254];
assign key[136]=and_result136[0]^and_result136[1]^and_result136[2]^and_result136[3]^and_result136[4]^and_result136[5]^and_result136[6]^and_result136[7]^and_result136[8]^and_result136[9]^and_result136[10]^and_result136[11]^and_result136[12]^and_result136[13]^and_result136[14]^and_result136[15]^and_result136[16]^and_result136[17]^and_result136[18]^and_result136[19]^and_result136[20]^and_result136[21]^and_result136[22]^and_result136[23]^and_result136[24]^and_result136[25]^and_result136[26]^and_result136[27]^and_result136[28]^and_result136[29]^and_result136[30]^and_result136[31]^and_result136[32]^and_result136[33]^and_result136[34]^and_result136[35]^and_result136[36]^and_result136[37]^and_result136[38]^and_result136[39]^and_result136[40]^and_result136[41]^and_result136[42]^and_result136[43]^and_result136[44]^and_result136[45]^and_result136[46]^and_result136[47]^and_result136[48]^and_result136[49]^and_result136[50]^and_result136[51]^and_result136[52]^and_result136[53]^and_result136[54]^and_result136[55]^and_result136[56]^and_result136[57]^and_result136[58]^and_result136[59]^and_result136[60]^and_result136[61]^and_result136[62]^and_result136[63]^and_result136[64]^and_result136[65]^and_result136[66]^and_result136[67]^and_result136[68]^and_result136[69]^and_result136[70]^and_result136[71]^and_result136[72]^and_result136[73]^and_result136[74]^and_result136[75]^and_result136[76]^and_result136[77]^and_result136[78]^and_result136[79]^and_result136[80]^and_result136[81]^and_result136[82]^and_result136[83]^and_result136[84]^and_result136[85]^and_result136[86]^and_result136[87]^and_result136[88]^and_result136[89]^and_result136[90]^and_result136[91]^and_result136[92]^and_result136[93]^and_result136[94]^and_result136[95]^and_result136[96]^and_result136[97]^and_result136[98]^and_result136[99]^and_result136[100]^and_result136[101]^and_result136[102]^and_result136[103]^and_result136[104]^and_result136[105]^and_result136[106]^and_result136[107]^and_result136[108]^and_result136[109]^and_result136[110]^and_result136[111]^and_result136[112]^and_result136[113]^and_result136[114]^and_result136[115]^and_result136[116]^and_result136[117]^and_result136[118]^and_result136[119]^and_result136[120]^and_result136[121]^and_result136[122]^and_result136[123]^and_result136[124]^and_result136[125]^and_result136[126]^and_result136[127]^and_result136[128]^and_result136[129]^and_result136[130]^and_result136[131]^and_result136[132]^and_result136[133]^and_result136[134]^and_result136[135]^and_result136[136]^and_result136[137]^and_result136[138]^and_result136[139]^and_result136[140]^and_result136[141]^and_result136[142]^and_result136[143]^and_result136[144]^and_result136[145]^and_result136[146]^and_result136[147]^and_result136[148]^and_result136[149]^and_result136[150]^and_result136[151]^and_result136[152]^and_result136[153]^and_result136[154]^and_result136[155]^and_result136[156]^and_result136[157]^and_result136[158]^and_result136[159]^and_result136[160]^and_result136[161]^and_result136[162]^and_result136[163]^and_result136[164]^and_result136[165]^and_result136[166]^and_result136[167]^and_result136[168]^and_result136[169]^and_result136[170]^and_result136[171]^and_result136[172]^and_result136[173]^and_result136[174]^and_result136[175]^and_result136[176]^and_result136[177]^and_result136[178]^and_result136[179]^and_result136[180]^and_result136[181]^and_result136[182]^and_result136[183]^and_result136[184]^and_result136[185]^and_result136[186]^and_result136[187]^and_result136[188]^and_result136[189]^and_result136[190]^and_result136[191]^and_result136[192]^and_result136[193]^and_result136[194]^and_result136[195]^and_result136[196]^and_result136[197]^and_result136[198]^and_result136[199]^and_result136[200]^and_result136[201]^and_result136[202]^and_result136[203]^and_result136[204]^and_result136[205]^and_result136[206]^and_result136[207]^and_result136[208]^and_result136[209]^and_result136[210]^and_result136[211]^and_result136[212]^and_result136[213]^and_result136[214]^and_result136[215]^and_result136[216]^and_result136[217]^and_result136[218]^and_result136[219]^and_result136[220]^and_result136[221]^and_result136[222]^and_result136[223]^and_result136[224]^and_result136[225]^and_result136[226]^and_result136[227]^and_result136[228]^and_result136[229]^and_result136[230]^and_result136[231]^and_result136[232]^and_result136[233]^and_result136[234]^and_result136[235]^and_result136[236]^and_result136[237]^and_result136[238]^and_result136[239]^and_result136[240]^and_result136[241]^and_result136[242]^and_result136[243]^and_result136[244]^and_result136[245]^and_result136[246]^and_result136[247]^and_result136[248]^and_result136[249]^and_result136[250]^and_result136[251]^and_result136[252]^and_result136[253]^and_result136[254];
assign key[137]=and_result137[0]^and_result137[1]^and_result137[2]^and_result137[3]^and_result137[4]^and_result137[5]^and_result137[6]^and_result137[7]^and_result137[8]^and_result137[9]^and_result137[10]^and_result137[11]^and_result137[12]^and_result137[13]^and_result137[14]^and_result137[15]^and_result137[16]^and_result137[17]^and_result137[18]^and_result137[19]^and_result137[20]^and_result137[21]^and_result137[22]^and_result137[23]^and_result137[24]^and_result137[25]^and_result137[26]^and_result137[27]^and_result137[28]^and_result137[29]^and_result137[30]^and_result137[31]^and_result137[32]^and_result137[33]^and_result137[34]^and_result137[35]^and_result137[36]^and_result137[37]^and_result137[38]^and_result137[39]^and_result137[40]^and_result137[41]^and_result137[42]^and_result137[43]^and_result137[44]^and_result137[45]^and_result137[46]^and_result137[47]^and_result137[48]^and_result137[49]^and_result137[50]^and_result137[51]^and_result137[52]^and_result137[53]^and_result137[54]^and_result137[55]^and_result137[56]^and_result137[57]^and_result137[58]^and_result137[59]^and_result137[60]^and_result137[61]^and_result137[62]^and_result137[63]^and_result137[64]^and_result137[65]^and_result137[66]^and_result137[67]^and_result137[68]^and_result137[69]^and_result137[70]^and_result137[71]^and_result137[72]^and_result137[73]^and_result137[74]^and_result137[75]^and_result137[76]^and_result137[77]^and_result137[78]^and_result137[79]^and_result137[80]^and_result137[81]^and_result137[82]^and_result137[83]^and_result137[84]^and_result137[85]^and_result137[86]^and_result137[87]^and_result137[88]^and_result137[89]^and_result137[90]^and_result137[91]^and_result137[92]^and_result137[93]^and_result137[94]^and_result137[95]^and_result137[96]^and_result137[97]^and_result137[98]^and_result137[99]^and_result137[100]^and_result137[101]^and_result137[102]^and_result137[103]^and_result137[104]^and_result137[105]^and_result137[106]^and_result137[107]^and_result137[108]^and_result137[109]^and_result137[110]^and_result137[111]^and_result137[112]^and_result137[113]^and_result137[114]^and_result137[115]^and_result137[116]^and_result137[117]^and_result137[118]^and_result137[119]^and_result137[120]^and_result137[121]^and_result137[122]^and_result137[123]^and_result137[124]^and_result137[125]^and_result137[126]^and_result137[127]^and_result137[128]^and_result137[129]^and_result137[130]^and_result137[131]^and_result137[132]^and_result137[133]^and_result137[134]^and_result137[135]^and_result137[136]^and_result137[137]^and_result137[138]^and_result137[139]^and_result137[140]^and_result137[141]^and_result137[142]^and_result137[143]^and_result137[144]^and_result137[145]^and_result137[146]^and_result137[147]^and_result137[148]^and_result137[149]^and_result137[150]^and_result137[151]^and_result137[152]^and_result137[153]^and_result137[154]^and_result137[155]^and_result137[156]^and_result137[157]^and_result137[158]^and_result137[159]^and_result137[160]^and_result137[161]^and_result137[162]^and_result137[163]^and_result137[164]^and_result137[165]^and_result137[166]^and_result137[167]^and_result137[168]^and_result137[169]^and_result137[170]^and_result137[171]^and_result137[172]^and_result137[173]^and_result137[174]^and_result137[175]^and_result137[176]^and_result137[177]^and_result137[178]^and_result137[179]^and_result137[180]^and_result137[181]^and_result137[182]^and_result137[183]^and_result137[184]^and_result137[185]^and_result137[186]^and_result137[187]^and_result137[188]^and_result137[189]^and_result137[190]^and_result137[191]^and_result137[192]^and_result137[193]^and_result137[194]^and_result137[195]^and_result137[196]^and_result137[197]^and_result137[198]^and_result137[199]^and_result137[200]^and_result137[201]^and_result137[202]^and_result137[203]^and_result137[204]^and_result137[205]^and_result137[206]^and_result137[207]^and_result137[208]^and_result137[209]^and_result137[210]^and_result137[211]^and_result137[212]^and_result137[213]^and_result137[214]^and_result137[215]^and_result137[216]^and_result137[217]^and_result137[218]^and_result137[219]^and_result137[220]^and_result137[221]^and_result137[222]^and_result137[223]^and_result137[224]^and_result137[225]^and_result137[226]^and_result137[227]^and_result137[228]^and_result137[229]^and_result137[230]^and_result137[231]^and_result137[232]^and_result137[233]^and_result137[234]^and_result137[235]^and_result137[236]^and_result137[237]^and_result137[238]^and_result137[239]^and_result137[240]^and_result137[241]^and_result137[242]^and_result137[243]^and_result137[244]^and_result137[245]^and_result137[246]^and_result137[247]^and_result137[248]^and_result137[249]^and_result137[250]^and_result137[251]^and_result137[252]^and_result137[253]^and_result137[254];
assign key[138]=and_result138[0]^and_result138[1]^and_result138[2]^and_result138[3]^and_result138[4]^and_result138[5]^and_result138[6]^and_result138[7]^and_result138[8]^and_result138[9]^and_result138[10]^and_result138[11]^and_result138[12]^and_result138[13]^and_result138[14]^and_result138[15]^and_result138[16]^and_result138[17]^and_result138[18]^and_result138[19]^and_result138[20]^and_result138[21]^and_result138[22]^and_result138[23]^and_result138[24]^and_result138[25]^and_result138[26]^and_result138[27]^and_result138[28]^and_result138[29]^and_result138[30]^and_result138[31]^and_result138[32]^and_result138[33]^and_result138[34]^and_result138[35]^and_result138[36]^and_result138[37]^and_result138[38]^and_result138[39]^and_result138[40]^and_result138[41]^and_result138[42]^and_result138[43]^and_result138[44]^and_result138[45]^and_result138[46]^and_result138[47]^and_result138[48]^and_result138[49]^and_result138[50]^and_result138[51]^and_result138[52]^and_result138[53]^and_result138[54]^and_result138[55]^and_result138[56]^and_result138[57]^and_result138[58]^and_result138[59]^and_result138[60]^and_result138[61]^and_result138[62]^and_result138[63]^and_result138[64]^and_result138[65]^and_result138[66]^and_result138[67]^and_result138[68]^and_result138[69]^and_result138[70]^and_result138[71]^and_result138[72]^and_result138[73]^and_result138[74]^and_result138[75]^and_result138[76]^and_result138[77]^and_result138[78]^and_result138[79]^and_result138[80]^and_result138[81]^and_result138[82]^and_result138[83]^and_result138[84]^and_result138[85]^and_result138[86]^and_result138[87]^and_result138[88]^and_result138[89]^and_result138[90]^and_result138[91]^and_result138[92]^and_result138[93]^and_result138[94]^and_result138[95]^and_result138[96]^and_result138[97]^and_result138[98]^and_result138[99]^and_result138[100]^and_result138[101]^and_result138[102]^and_result138[103]^and_result138[104]^and_result138[105]^and_result138[106]^and_result138[107]^and_result138[108]^and_result138[109]^and_result138[110]^and_result138[111]^and_result138[112]^and_result138[113]^and_result138[114]^and_result138[115]^and_result138[116]^and_result138[117]^and_result138[118]^and_result138[119]^and_result138[120]^and_result138[121]^and_result138[122]^and_result138[123]^and_result138[124]^and_result138[125]^and_result138[126]^and_result138[127]^and_result138[128]^and_result138[129]^and_result138[130]^and_result138[131]^and_result138[132]^and_result138[133]^and_result138[134]^and_result138[135]^and_result138[136]^and_result138[137]^and_result138[138]^and_result138[139]^and_result138[140]^and_result138[141]^and_result138[142]^and_result138[143]^and_result138[144]^and_result138[145]^and_result138[146]^and_result138[147]^and_result138[148]^and_result138[149]^and_result138[150]^and_result138[151]^and_result138[152]^and_result138[153]^and_result138[154]^and_result138[155]^and_result138[156]^and_result138[157]^and_result138[158]^and_result138[159]^and_result138[160]^and_result138[161]^and_result138[162]^and_result138[163]^and_result138[164]^and_result138[165]^and_result138[166]^and_result138[167]^and_result138[168]^and_result138[169]^and_result138[170]^and_result138[171]^and_result138[172]^and_result138[173]^and_result138[174]^and_result138[175]^and_result138[176]^and_result138[177]^and_result138[178]^and_result138[179]^and_result138[180]^and_result138[181]^and_result138[182]^and_result138[183]^and_result138[184]^and_result138[185]^and_result138[186]^and_result138[187]^and_result138[188]^and_result138[189]^and_result138[190]^and_result138[191]^and_result138[192]^and_result138[193]^and_result138[194]^and_result138[195]^and_result138[196]^and_result138[197]^and_result138[198]^and_result138[199]^and_result138[200]^and_result138[201]^and_result138[202]^and_result138[203]^and_result138[204]^and_result138[205]^and_result138[206]^and_result138[207]^and_result138[208]^and_result138[209]^and_result138[210]^and_result138[211]^and_result138[212]^and_result138[213]^and_result138[214]^and_result138[215]^and_result138[216]^and_result138[217]^and_result138[218]^and_result138[219]^and_result138[220]^and_result138[221]^and_result138[222]^and_result138[223]^and_result138[224]^and_result138[225]^and_result138[226]^and_result138[227]^and_result138[228]^and_result138[229]^and_result138[230]^and_result138[231]^and_result138[232]^and_result138[233]^and_result138[234]^and_result138[235]^and_result138[236]^and_result138[237]^and_result138[238]^and_result138[239]^and_result138[240]^and_result138[241]^and_result138[242]^and_result138[243]^and_result138[244]^and_result138[245]^and_result138[246]^and_result138[247]^and_result138[248]^and_result138[249]^and_result138[250]^and_result138[251]^and_result138[252]^and_result138[253]^and_result138[254];
assign key[139]=and_result139[0]^and_result139[1]^and_result139[2]^and_result139[3]^and_result139[4]^and_result139[5]^and_result139[6]^and_result139[7]^and_result139[8]^and_result139[9]^and_result139[10]^and_result139[11]^and_result139[12]^and_result139[13]^and_result139[14]^and_result139[15]^and_result139[16]^and_result139[17]^and_result139[18]^and_result139[19]^and_result139[20]^and_result139[21]^and_result139[22]^and_result139[23]^and_result139[24]^and_result139[25]^and_result139[26]^and_result139[27]^and_result139[28]^and_result139[29]^and_result139[30]^and_result139[31]^and_result139[32]^and_result139[33]^and_result139[34]^and_result139[35]^and_result139[36]^and_result139[37]^and_result139[38]^and_result139[39]^and_result139[40]^and_result139[41]^and_result139[42]^and_result139[43]^and_result139[44]^and_result139[45]^and_result139[46]^and_result139[47]^and_result139[48]^and_result139[49]^and_result139[50]^and_result139[51]^and_result139[52]^and_result139[53]^and_result139[54]^and_result139[55]^and_result139[56]^and_result139[57]^and_result139[58]^and_result139[59]^and_result139[60]^and_result139[61]^and_result139[62]^and_result139[63]^and_result139[64]^and_result139[65]^and_result139[66]^and_result139[67]^and_result139[68]^and_result139[69]^and_result139[70]^and_result139[71]^and_result139[72]^and_result139[73]^and_result139[74]^and_result139[75]^and_result139[76]^and_result139[77]^and_result139[78]^and_result139[79]^and_result139[80]^and_result139[81]^and_result139[82]^and_result139[83]^and_result139[84]^and_result139[85]^and_result139[86]^and_result139[87]^and_result139[88]^and_result139[89]^and_result139[90]^and_result139[91]^and_result139[92]^and_result139[93]^and_result139[94]^and_result139[95]^and_result139[96]^and_result139[97]^and_result139[98]^and_result139[99]^and_result139[100]^and_result139[101]^and_result139[102]^and_result139[103]^and_result139[104]^and_result139[105]^and_result139[106]^and_result139[107]^and_result139[108]^and_result139[109]^and_result139[110]^and_result139[111]^and_result139[112]^and_result139[113]^and_result139[114]^and_result139[115]^and_result139[116]^and_result139[117]^and_result139[118]^and_result139[119]^and_result139[120]^and_result139[121]^and_result139[122]^and_result139[123]^and_result139[124]^and_result139[125]^and_result139[126]^and_result139[127]^and_result139[128]^and_result139[129]^and_result139[130]^and_result139[131]^and_result139[132]^and_result139[133]^and_result139[134]^and_result139[135]^and_result139[136]^and_result139[137]^and_result139[138]^and_result139[139]^and_result139[140]^and_result139[141]^and_result139[142]^and_result139[143]^and_result139[144]^and_result139[145]^and_result139[146]^and_result139[147]^and_result139[148]^and_result139[149]^and_result139[150]^and_result139[151]^and_result139[152]^and_result139[153]^and_result139[154]^and_result139[155]^and_result139[156]^and_result139[157]^and_result139[158]^and_result139[159]^and_result139[160]^and_result139[161]^and_result139[162]^and_result139[163]^and_result139[164]^and_result139[165]^and_result139[166]^and_result139[167]^and_result139[168]^and_result139[169]^and_result139[170]^and_result139[171]^and_result139[172]^and_result139[173]^and_result139[174]^and_result139[175]^and_result139[176]^and_result139[177]^and_result139[178]^and_result139[179]^and_result139[180]^and_result139[181]^and_result139[182]^and_result139[183]^and_result139[184]^and_result139[185]^and_result139[186]^and_result139[187]^and_result139[188]^and_result139[189]^and_result139[190]^and_result139[191]^and_result139[192]^and_result139[193]^and_result139[194]^and_result139[195]^and_result139[196]^and_result139[197]^and_result139[198]^and_result139[199]^and_result139[200]^and_result139[201]^and_result139[202]^and_result139[203]^and_result139[204]^and_result139[205]^and_result139[206]^and_result139[207]^and_result139[208]^and_result139[209]^and_result139[210]^and_result139[211]^and_result139[212]^and_result139[213]^and_result139[214]^and_result139[215]^and_result139[216]^and_result139[217]^and_result139[218]^and_result139[219]^and_result139[220]^and_result139[221]^and_result139[222]^and_result139[223]^and_result139[224]^and_result139[225]^and_result139[226]^and_result139[227]^and_result139[228]^and_result139[229]^and_result139[230]^and_result139[231]^and_result139[232]^and_result139[233]^and_result139[234]^and_result139[235]^and_result139[236]^and_result139[237]^and_result139[238]^and_result139[239]^and_result139[240]^and_result139[241]^and_result139[242]^and_result139[243]^and_result139[244]^and_result139[245]^and_result139[246]^and_result139[247]^and_result139[248]^and_result139[249]^and_result139[250]^and_result139[251]^and_result139[252]^and_result139[253]^and_result139[254];
assign key[140]=and_result140[0]^and_result140[1]^and_result140[2]^and_result140[3]^and_result140[4]^and_result140[5]^and_result140[6]^and_result140[7]^and_result140[8]^and_result140[9]^and_result140[10]^and_result140[11]^and_result140[12]^and_result140[13]^and_result140[14]^and_result140[15]^and_result140[16]^and_result140[17]^and_result140[18]^and_result140[19]^and_result140[20]^and_result140[21]^and_result140[22]^and_result140[23]^and_result140[24]^and_result140[25]^and_result140[26]^and_result140[27]^and_result140[28]^and_result140[29]^and_result140[30]^and_result140[31]^and_result140[32]^and_result140[33]^and_result140[34]^and_result140[35]^and_result140[36]^and_result140[37]^and_result140[38]^and_result140[39]^and_result140[40]^and_result140[41]^and_result140[42]^and_result140[43]^and_result140[44]^and_result140[45]^and_result140[46]^and_result140[47]^and_result140[48]^and_result140[49]^and_result140[50]^and_result140[51]^and_result140[52]^and_result140[53]^and_result140[54]^and_result140[55]^and_result140[56]^and_result140[57]^and_result140[58]^and_result140[59]^and_result140[60]^and_result140[61]^and_result140[62]^and_result140[63]^and_result140[64]^and_result140[65]^and_result140[66]^and_result140[67]^and_result140[68]^and_result140[69]^and_result140[70]^and_result140[71]^and_result140[72]^and_result140[73]^and_result140[74]^and_result140[75]^and_result140[76]^and_result140[77]^and_result140[78]^and_result140[79]^and_result140[80]^and_result140[81]^and_result140[82]^and_result140[83]^and_result140[84]^and_result140[85]^and_result140[86]^and_result140[87]^and_result140[88]^and_result140[89]^and_result140[90]^and_result140[91]^and_result140[92]^and_result140[93]^and_result140[94]^and_result140[95]^and_result140[96]^and_result140[97]^and_result140[98]^and_result140[99]^and_result140[100]^and_result140[101]^and_result140[102]^and_result140[103]^and_result140[104]^and_result140[105]^and_result140[106]^and_result140[107]^and_result140[108]^and_result140[109]^and_result140[110]^and_result140[111]^and_result140[112]^and_result140[113]^and_result140[114]^and_result140[115]^and_result140[116]^and_result140[117]^and_result140[118]^and_result140[119]^and_result140[120]^and_result140[121]^and_result140[122]^and_result140[123]^and_result140[124]^and_result140[125]^and_result140[126]^and_result140[127]^and_result140[128]^and_result140[129]^and_result140[130]^and_result140[131]^and_result140[132]^and_result140[133]^and_result140[134]^and_result140[135]^and_result140[136]^and_result140[137]^and_result140[138]^and_result140[139]^and_result140[140]^and_result140[141]^and_result140[142]^and_result140[143]^and_result140[144]^and_result140[145]^and_result140[146]^and_result140[147]^and_result140[148]^and_result140[149]^and_result140[150]^and_result140[151]^and_result140[152]^and_result140[153]^and_result140[154]^and_result140[155]^and_result140[156]^and_result140[157]^and_result140[158]^and_result140[159]^and_result140[160]^and_result140[161]^and_result140[162]^and_result140[163]^and_result140[164]^and_result140[165]^and_result140[166]^and_result140[167]^and_result140[168]^and_result140[169]^and_result140[170]^and_result140[171]^and_result140[172]^and_result140[173]^and_result140[174]^and_result140[175]^and_result140[176]^and_result140[177]^and_result140[178]^and_result140[179]^and_result140[180]^and_result140[181]^and_result140[182]^and_result140[183]^and_result140[184]^and_result140[185]^and_result140[186]^and_result140[187]^and_result140[188]^and_result140[189]^and_result140[190]^and_result140[191]^and_result140[192]^and_result140[193]^and_result140[194]^and_result140[195]^and_result140[196]^and_result140[197]^and_result140[198]^and_result140[199]^and_result140[200]^and_result140[201]^and_result140[202]^and_result140[203]^and_result140[204]^and_result140[205]^and_result140[206]^and_result140[207]^and_result140[208]^and_result140[209]^and_result140[210]^and_result140[211]^and_result140[212]^and_result140[213]^and_result140[214]^and_result140[215]^and_result140[216]^and_result140[217]^and_result140[218]^and_result140[219]^and_result140[220]^and_result140[221]^and_result140[222]^and_result140[223]^and_result140[224]^and_result140[225]^and_result140[226]^and_result140[227]^and_result140[228]^and_result140[229]^and_result140[230]^and_result140[231]^and_result140[232]^and_result140[233]^and_result140[234]^and_result140[235]^and_result140[236]^and_result140[237]^and_result140[238]^and_result140[239]^and_result140[240]^and_result140[241]^and_result140[242]^and_result140[243]^and_result140[244]^and_result140[245]^and_result140[246]^and_result140[247]^and_result140[248]^and_result140[249]^and_result140[250]^and_result140[251]^and_result140[252]^and_result140[253]^and_result140[254];
assign key[141]=and_result141[0]^and_result141[1]^and_result141[2]^and_result141[3]^and_result141[4]^and_result141[5]^and_result141[6]^and_result141[7]^and_result141[8]^and_result141[9]^and_result141[10]^and_result141[11]^and_result141[12]^and_result141[13]^and_result141[14]^and_result141[15]^and_result141[16]^and_result141[17]^and_result141[18]^and_result141[19]^and_result141[20]^and_result141[21]^and_result141[22]^and_result141[23]^and_result141[24]^and_result141[25]^and_result141[26]^and_result141[27]^and_result141[28]^and_result141[29]^and_result141[30]^and_result141[31]^and_result141[32]^and_result141[33]^and_result141[34]^and_result141[35]^and_result141[36]^and_result141[37]^and_result141[38]^and_result141[39]^and_result141[40]^and_result141[41]^and_result141[42]^and_result141[43]^and_result141[44]^and_result141[45]^and_result141[46]^and_result141[47]^and_result141[48]^and_result141[49]^and_result141[50]^and_result141[51]^and_result141[52]^and_result141[53]^and_result141[54]^and_result141[55]^and_result141[56]^and_result141[57]^and_result141[58]^and_result141[59]^and_result141[60]^and_result141[61]^and_result141[62]^and_result141[63]^and_result141[64]^and_result141[65]^and_result141[66]^and_result141[67]^and_result141[68]^and_result141[69]^and_result141[70]^and_result141[71]^and_result141[72]^and_result141[73]^and_result141[74]^and_result141[75]^and_result141[76]^and_result141[77]^and_result141[78]^and_result141[79]^and_result141[80]^and_result141[81]^and_result141[82]^and_result141[83]^and_result141[84]^and_result141[85]^and_result141[86]^and_result141[87]^and_result141[88]^and_result141[89]^and_result141[90]^and_result141[91]^and_result141[92]^and_result141[93]^and_result141[94]^and_result141[95]^and_result141[96]^and_result141[97]^and_result141[98]^and_result141[99]^and_result141[100]^and_result141[101]^and_result141[102]^and_result141[103]^and_result141[104]^and_result141[105]^and_result141[106]^and_result141[107]^and_result141[108]^and_result141[109]^and_result141[110]^and_result141[111]^and_result141[112]^and_result141[113]^and_result141[114]^and_result141[115]^and_result141[116]^and_result141[117]^and_result141[118]^and_result141[119]^and_result141[120]^and_result141[121]^and_result141[122]^and_result141[123]^and_result141[124]^and_result141[125]^and_result141[126]^and_result141[127]^and_result141[128]^and_result141[129]^and_result141[130]^and_result141[131]^and_result141[132]^and_result141[133]^and_result141[134]^and_result141[135]^and_result141[136]^and_result141[137]^and_result141[138]^and_result141[139]^and_result141[140]^and_result141[141]^and_result141[142]^and_result141[143]^and_result141[144]^and_result141[145]^and_result141[146]^and_result141[147]^and_result141[148]^and_result141[149]^and_result141[150]^and_result141[151]^and_result141[152]^and_result141[153]^and_result141[154]^and_result141[155]^and_result141[156]^and_result141[157]^and_result141[158]^and_result141[159]^and_result141[160]^and_result141[161]^and_result141[162]^and_result141[163]^and_result141[164]^and_result141[165]^and_result141[166]^and_result141[167]^and_result141[168]^and_result141[169]^and_result141[170]^and_result141[171]^and_result141[172]^and_result141[173]^and_result141[174]^and_result141[175]^and_result141[176]^and_result141[177]^and_result141[178]^and_result141[179]^and_result141[180]^and_result141[181]^and_result141[182]^and_result141[183]^and_result141[184]^and_result141[185]^and_result141[186]^and_result141[187]^and_result141[188]^and_result141[189]^and_result141[190]^and_result141[191]^and_result141[192]^and_result141[193]^and_result141[194]^and_result141[195]^and_result141[196]^and_result141[197]^and_result141[198]^and_result141[199]^and_result141[200]^and_result141[201]^and_result141[202]^and_result141[203]^and_result141[204]^and_result141[205]^and_result141[206]^and_result141[207]^and_result141[208]^and_result141[209]^and_result141[210]^and_result141[211]^and_result141[212]^and_result141[213]^and_result141[214]^and_result141[215]^and_result141[216]^and_result141[217]^and_result141[218]^and_result141[219]^and_result141[220]^and_result141[221]^and_result141[222]^and_result141[223]^and_result141[224]^and_result141[225]^and_result141[226]^and_result141[227]^and_result141[228]^and_result141[229]^and_result141[230]^and_result141[231]^and_result141[232]^and_result141[233]^and_result141[234]^and_result141[235]^and_result141[236]^and_result141[237]^and_result141[238]^and_result141[239]^and_result141[240]^and_result141[241]^and_result141[242]^and_result141[243]^and_result141[244]^and_result141[245]^and_result141[246]^and_result141[247]^and_result141[248]^and_result141[249]^and_result141[250]^and_result141[251]^and_result141[252]^and_result141[253]^and_result141[254];
assign key[142]=and_result142[0]^and_result142[1]^and_result142[2]^and_result142[3]^and_result142[4]^and_result142[5]^and_result142[6]^and_result142[7]^and_result142[8]^and_result142[9]^and_result142[10]^and_result142[11]^and_result142[12]^and_result142[13]^and_result142[14]^and_result142[15]^and_result142[16]^and_result142[17]^and_result142[18]^and_result142[19]^and_result142[20]^and_result142[21]^and_result142[22]^and_result142[23]^and_result142[24]^and_result142[25]^and_result142[26]^and_result142[27]^and_result142[28]^and_result142[29]^and_result142[30]^and_result142[31]^and_result142[32]^and_result142[33]^and_result142[34]^and_result142[35]^and_result142[36]^and_result142[37]^and_result142[38]^and_result142[39]^and_result142[40]^and_result142[41]^and_result142[42]^and_result142[43]^and_result142[44]^and_result142[45]^and_result142[46]^and_result142[47]^and_result142[48]^and_result142[49]^and_result142[50]^and_result142[51]^and_result142[52]^and_result142[53]^and_result142[54]^and_result142[55]^and_result142[56]^and_result142[57]^and_result142[58]^and_result142[59]^and_result142[60]^and_result142[61]^and_result142[62]^and_result142[63]^and_result142[64]^and_result142[65]^and_result142[66]^and_result142[67]^and_result142[68]^and_result142[69]^and_result142[70]^and_result142[71]^and_result142[72]^and_result142[73]^and_result142[74]^and_result142[75]^and_result142[76]^and_result142[77]^and_result142[78]^and_result142[79]^and_result142[80]^and_result142[81]^and_result142[82]^and_result142[83]^and_result142[84]^and_result142[85]^and_result142[86]^and_result142[87]^and_result142[88]^and_result142[89]^and_result142[90]^and_result142[91]^and_result142[92]^and_result142[93]^and_result142[94]^and_result142[95]^and_result142[96]^and_result142[97]^and_result142[98]^and_result142[99]^and_result142[100]^and_result142[101]^and_result142[102]^and_result142[103]^and_result142[104]^and_result142[105]^and_result142[106]^and_result142[107]^and_result142[108]^and_result142[109]^and_result142[110]^and_result142[111]^and_result142[112]^and_result142[113]^and_result142[114]^and_result142[115]^and_result142[116]^and_result142[117]^and_result142[118]^and_result142[119]^and_result142[120]^and_result142[121]^and_result142[122]^and_result142[123]^and_result142[124]^and_result142[125]^and_result142[126]^and_result142[127]^and_result142[128]^and_result142[129]^and_result142[130]^and_result142[131]^and_result142[132]^and_result142[133]^and_result142[134]^and_result142[135]^and_result142[136]^and_result142[137]^and_result142[138]^and_result142[139]^and_result142[140]^and_result142[141]^and_result142[142]^and_result142[143]^and_result142[144]^and_result142[145]^and_result142[146]^and_result142[147]^and_result142[148]^and_result142[149]^and_result142[150]^and_result142[151]^and_result142[152]^and_result142[153]^and_result142[154]^and_result142[155]^and_result142[156]^and_result142[157]^and_result142[158]^and_result142[159]^and_result142[160]^and_result142[161]^and_result142[162]^and_result142[163]^and_result142[164]^and_result142[165]^and_result142[166]^and_result142[167]^and_result142[168]^and_result142[169]^and_result142[170]^and_result142[171]^and_result142[172]^and_result142[173]^and_result142[174]^and_result142[175]^and_result142[176]^and_result142[177]^and_result142[178]^and_result142[179]^and_result142[180]^and_result142[181]^and_result142[182]^and_result142[183]^and_result142[184]^and_result142[185]^and_result142[186]^and_result142[187]^and_result142[188]^and_result142[189]^and_result142[190]^and_result142[191]^and_result142[192]^and_result142[193]^and_result142[194]^and_result142[195]^and_result142[196]^and_result142[197]^and_result142[198]^and_result142[199]^and_result142[200]^and_result142[201]^and_result142[202]^and_result142[203]^and_result142[204]^and_result142[205]^and_result142[206]^and_result142[207]^and_result142[208]^and_result142[209]^and_result142[210]^and_result142[211]^and_result142[212]^and_result142[213]^and_result142[214]^and_result142[215]^and_result142[216]^and_result142[217]^and_result142[218]^and_result142[219]^and_result142[220]^and_result142[221]^and_result142[222]^and_result142[223]^and_result142[224]^and_result142[225]^and_result142[226]^and_result142[227]^and_result142[228]^and_result142[229]^and_result142[230]^and_result142[231]^and_result142[232]^and_result142[233]^and_result142[234]^and_result142[235]^and_result142[236]^and_result142[237]^and_result142[238]^and_result142[239]^and_result142[240]^and_result142[241]^and_result142[242]^and_result142[243]^and_result142[244]^and_result142[245]^and_result142[246]^and_result142[247]^and_result142[248]^and_result142[249]^and_result142[250]^and_result142[251]^and_result142[252]^and_result142[253]^and_result142[254];
assign key[143]=and_result143[0]^and_result143[1]^and_result143[2]^and_result143[3]^and_result143[4]^and_result143[5]^and_result143[6]^and_result143[7]^and_result143[8]^and_result143[9]^and_result143[10]^and_result143[11]^and_result143[12]^and_result143[13]^and_result143[14]^and_result143[15]^and_result143[16]^and_result143[17]^and_result143[18]^and_result143[19]^and_result143[20]^and_result143[21]^and_result143[22]^and_result143[23]^and_result143[24]^and_result143[25]^and_result143[26]^and_result143[27]^and_result143[28]^and_result143[29]^and_result143[30]^and_result143[31]^and_result143[32]^and_result143[33]^and_result143[34]^and_result143[35]^and_result143[36]^and_result143[37]^and_result143[38]^and_result143[39]^and_result143[40]^and_result143[41]^and_result143[42]^and_result143[43]^and_result143[44]^and_result143[45]^and_result143[46]^and_result143[47]^and_result143[48]^and_result143[49]^and_result143[50]^and_result143[51]^and_result143[52]^and_result143[53]^and_result143[54]^and_result143[55]^and_result143[56]^and_result143[57]^and_result143[58]^and_result143[59]^and_result143[60]^and_result143[61]^and_result143[62]^and_result143[63]^and_result143[64]^and_result143[65]^and_result143[66]^and_result143[67]^and_result143[68]^and_result143[69]^and_result143[70]^and_result143[71]^and_result143[72]^and_result143[73]^and_result143[74]^and_result143[75]^and_result143[76]^and_result143[77]^and_result143[78]^and_result143[79]^and_result143[80]^and_result143[81]^and_result143[82]^and_result143[83]^and_result143[84]^and_result143[85]^and_result143[86]^and_result143[87]^and_result143[88]^and_result143[89]^and_result143[90]^and_result143[91]^and_result143[92]^and_result143[93]^and_result143[94]^and_result143[95]^and_result143[96]^and_result143[97]^and_result143[98]^and_result143[99]^and_result143[100]^and_result143[101]^and_result143[102]^and_result143[103]^and_result143[104]^and_result143[105]^and_result143[106]^and_result143[107]^and_result143[108]^and_result143[109]^and_result143[110]^and_result143[111]^and_result143[112]^and_result143[113]^and_result143[114]^and_result143[115]^and_result143[116]^and_result143[117]^and_result143[118]^and_result143[119]^and_result143[120]^and_result143[121]^and_result143[122]^and_result143[123]^and_result143[124]^and_result143[125]^and_result143[126]^and_result143[127]^and_result143[128]^and_result143[129]^and_result143[130]^and_result143[131]^and_result143[132]^and_result143[133]^and_result143[134]^and_result143[135]^and_result143[136]^and_result143[137]^and_result143[138]^and_result143[139]^and_result143[140]^and_result143[141]^and_result143[142]^and_result143[143]^and_result143[144]^and_result143[145]^and_result143[146]^and_result143[147]^and_result143[148]^and_result143[149]^and_result143[150]^and_result143[151]^and_result143[152]^and_result143[153]^and_result143[154]^and_result143[155]^and_result143[156]^and_result143[157]^and_result143[158]^and_result143[159]^and_result143[160]^and_result143[161]^and_result143[162]^and_result143[163]^and_result143[164]^and_result143[165]^and_result143[166]^and_result143[167]^and_result143[168]^and_result143[169]^and_result143[170]^and_result143[171]^and_result143[172]^and_result143[173]^and_result143[174]^and_result143[175]^and_result143[176]^and_result143[177]^and_result143[178]^and_result143[179]^and_result143[180]^and_result143[181]^and_result143[182]^and_result143[183]^and_result143[184]^and_result143[185]^and_result143[186]^and_result143[187]^and_result143[188]^and_result143[189]^and_result143[190]^and_result143[191]^and_result143[192]^and_result143[193]^and_result143[194]^and_result143[195]^and_result143[196]^and_result143[197]^and_result143[198]^and_result143[199]^and_result143[200]^and_result143[201]^and_result143[202]^and_result143[203]^and_result143[204]^and_result143[205]^and_result143[206]^and_result143[207]^and_result143[208]^and_result143[209]^and_result143[210]^and_result143[211]^and_result143[212]^and_result143[213]^and_result143[214]^and_result143[215]^and_result143[216]^and_result143[217]^and_result143[218]^and_result143[219]^and_result143[220]^and_result143[221]^and_result143[222]^and_result143[223]^and_result143[224]^and_result143[225]^and_result143[226]^and_result143[227]^and_result143[228]^and_result143[229]^and_result143[230]^and_result143[231]^and_result143[232]^and_result143[233]^and_result143[234]^and_result143[235]^and_result143[236]^and_result143[237]^and_result143[238]^and_result143[239]^and_result143[240]^and_result143[241]^and_result143[242]^and_result143[243]^and_result143[244]^and_result143[245]^and_result143[246]^and_result143[247]^and_result143[248]^and_result143[249]^and_result143[250]^and_result143[251]^and_result143[252]^and_result143[253]^and_result143[254];
assign key[144]=and_result144[0]^and_result144[1]^and_result144[2]^and_result144[3]^and_result144[4]^and_result144[5]^and_result144[6]^and_result144[7]^and_result144[8]^and_result144[9]^and_result144[10]^and_result144[11]^and_result144[12]^and_result144[13]^and_result144[14]^and_result144[15]^and_result144[16]^and_result144[17]^and_result144[18]^and_result144[19]^and_result144[20]^and_result144[21]^and_result144[22]^and_result144[23]^and_result144[24]^and_result144[25]^and_result144[26]^and_result144[27]^and_result144[28]^and_result144[29]^and_result144[30]^and_result144[31]^and_result144[32]^and_result144[33]^and_result144[34]^and_result144[35]^and_result144[36]^and_result144[37]^and_result144[38]^and_result144[39]^and_result144[40]^and_result144[41]^and_result144[42]^and_result144[43]^and_result144[44]^and_result144[45]^and_result144[46]^and_result144[47]^and_result144[48]^and_result144[49]^and_result144[50]^and_result144[51]^and_result144[52]^and_result144[53]^and_result144[54]^and_result144[55]^and_result144[56]^and_result144[57]^and_result144[58]^and_result144[59]^and_result144[60]^and_result144[61]^and_result144[62]^and_result144[63]^and_result144[64]^and_result144[65]^and_result144[66]^and_result144[67]^and_result144[68]^and_result144[69]^and_result144[70]^and_result144[71]^and_result144[72]^and_result144[73]^and_result144[74]^and_result144[75]^and_result144[76]^and_result144[77]^and_result144[78]^and_result144[79]^and_result144[80]^and_result144[81]^and_result144[82]^and_result144[83]^and_result144[84]^and_result144[85]^and_result144[86]^and_result144[87]^and_result144[88]^and_result144[89]^and_result144[90]^and_result144[91]^and_result144[92]^and_result144[93]^and_result144[94]^and_result144[95]^and_result144[96]^and_result144[97]^and_result144[98]^and_result144[99]^and_result144[100]^and_result144[101]^and_result144[102]^and_result144[103]^and_result144[104]^and_result144[105]^and_result144[106]^and_result144[107]^and_result144[108]^and_result144[109]^and_result144[110]^and_result144[111]^and_result144[112]^and_result144[113]^and_result144[114]^and_result144[115]^and_result144[116]^and_result144[117]^and_result144[118]^and_result144[119]^and_result144[120]^and_result144[121]^and_result144[122]^and_result144[123]^and_result144[124]^and_result144[125]^and_result144[126]^and_result144[127]^and_result144[128]^and_result144[129]^and_result144[130]^and_result144[131]^and_result144[132]^and_result144[133]^and_result144[134]^and_result144[135]^and_result144[136]^and_result144[137]^and_result144[138]^and_result144[139]^and_result144[140]^and_result144[141]^and_result144[142]^and_result144[143]^and_result144[144]^and_result144[145]^and_result144[146]^and_result144[147]^and_result144[148]^and_result144[149]^and_result144[150]^and_result144[151]^and_result144[152]^and_result144[153]^and_result144[154]^and_result144[155]^and_result144[156]^and_result144[157]^and_result144[158]^and_result144[159]^and_result144[160]^and_result144[161]^and_result144[162]^and_result144[163]^and_result144[164]^and_result144[165]^and_result144[166]^and_result144[167]^and_result144[168]^and_result144[169]^and_result144[170]^and_result144[171]^and_result144[172]^and_result144[173]^and_result144[174]^and_result144[175]^and_result144[176]^and_result144[177]^and_result144[178]^and_result144[179]^and_result144[180]^and_result144[181]^and_result144[182]^and_result144[183]^and_result144[184]^and_result144[185]^and_result144[186]^and_result144[187]^and_result144[188]^and_result144[189]^and_result144[190]^and_result144[191]^and_result144[192]^and_result144[193]^and_result144[194]^and_result144[195]^and_result144[196]^and_result144[197]^and_result144[198]^and_result144[199]^and_result144[200]^and_result144[201]^and_result144[202]^and_result144[203]^and_result144[204]^and_result144[205]^and_result144[206]^and_result144[207]^and_result144[208]^and_result144[209]^and_result144[210]^and_result144[211]^and_result144[212]^and_result144[213]^and_result144[214]^and_result144[215]^and_result144[216]^and_result144[217]^and_result144[218]^and_result144[219]^and_result144[220]^and_result144[221]^and_result144[222]^and_result144[223]^and_result144[224]^and_result144[225]^and_result144[226]^and_result144[227]^and_result144[228]^and_result144[229]^and_result144[230]^and_result144[231]^and_result144[232]^and_result144[233]^and_result144[234]^and_result144[235]^and_result144[236]^and_result144[237]^and_result144[238]^and_result144[239]^and_result144[240]^and_result144[241]^and_result144[242]^and_result144[243]^and_result144[244]^and_result144[245]^and_result144[246]^and_result144[247]^and_result144[248]^and_result144[249]^and_result144[250]^and_result144[251]^and_result144[252]^and_result144[253]^and_result144[254];
assign key[145]=and_result145[0]^and_result145[1]^and_result145[2]^and_result145[3]^and_result145[4]^and_result145[5]^and_result145[6]^and_result145[7]^and_result145[8]^and_result145[9]^and_result145[10]^and_result145[11]^and_result145[12]^and_result145[13]^and_result145[14]^and_result145[15]^and_result145[16]^and_result145[17]^and_result145[18]^and_result145[19]^and_result145[20]^and_result145[21]^and_result145[22]^and_result145[23]^and_result145[24]^and_result145[25]^and_result145[26]^and_result145[27]^and_result145[28]^and_result145[29]^and_result145[30]^and_result145[31]^and_result145[32]^and_result145[33]^and_result145[34]^and_result145[35]^and_result145[36]^and_result145[37]^and_result145[38]^and_result145[39]^and_result145[40]^and_result145[41]^and_result145[42]^and_result145[43]^and_result145[44]^and_result145[45]^and_result145[46]^and_result145[47]^and_result145[48]^and_result145[49]^and_result145[50]^and_result145[51]^and_result145[52]^and_result145[53]^and_result145[54]^and_result145[55]^and_result145[56]^and_result145[57]^and_result145[58]^and_result145[59]^and_result145[60]^and_result145[61]^and_result145[62]^and_result145[63]^and_result145[64]^and_result145[65]^and_result145[66]^and_result145[67]^and_result145[68]^and_result145[69]^and_result145[70]^and_result145[71]^and_result145[72]^and_result145[73]^and_result145[74]^and_result145[75]^and_result145[76]^and_result145[77]^and_result145[78]^and_result145[79]^and_result145[80]^and_result145[81]^and_result145[82]^and_result145[83]^and_result145[84]^and_result145[85]^and_result145[86]^and_result145[87]^and_result145[88]^and_result145[89]^and_result145[90]^and_result145[91]^and_result145[92]^and_result145[93]^and_result145[94]^and_result145[95]^and_result145[96]^and_result145[97]^and_result145[98]^and_result145[99]^and_result145[100]^and_result145[101]^and_result145[102]^and_result145[103]^and_result145[104]^and_result145[105]^and_result145[106]^and_result145[107]^and_result145[108]^and_result145[109]^and_result145[110]^and_result145[111]^and_result145[112]^and_result145[113]^and_result145[114]^and_result145[115]^and_result145[116]^and_result145[117]^and_result145[118]^and_result145[119]^and_result145[120]^and_result145[121]^and_result145[122]^and_result145[123]^and_result145[124]^and_result145[125]^and_result145[126]^and_result145[127]^and_result145[128]^and_result145[129]^and_result145[130]^and_result145[131]^and_result145[132]^and_result145[133]^and_result145[134]^and_result145[135]^and_result145[136]^and_result145[137]^and_result145[138]^and_result145[139]^and_result145[140]^and_result145[141]^and_result145[142]^and_result145[143]^and_result145[144]^and_result145[145]^and_result145[146]^and_result145[147]^and_result145[148]^and_result145[149]^and_result145[150]^and_result145[151]^and_result145[152]^and_result145[153]^and_result145[154]^and_result145[155]^and_result145[156]^and_result145[157]^and_result145[158]^and_result145[159]^and_result145[160]^and_result145[161]^and_result145[162]^and_result145[163]^and_result145[164]^and_result145[165]^and_result145[166]^and_result145[167]^and_result145[168]^and_result145[169]^and_result145[170]^and_result145[171]^and_result145[172]^and_result145[173]^and_result145[174]^and_result145[175]^and_result145[176]^and_result145[177]^and_result145[178]^and_result145[179]^and_result145[180]^and_result145[181]^and_result145[182]^and_result145[183]^and_result145[184]^and_result145[185]^and_result145[186]^and_result145[187]^and_result145[188]^and_result145[189]^and_result145[190]^and_result145[191]^and_result145[192]^and_result145[193]^and_result145[194]^and_result145[195]^and_result145[196]^and_result145[197]^and_result145[198]^and_result145[199]^and_result145[200]^and_result145[201]^and_result145[202]^and_result145[203]^and_result145[204]^and_result145[205]^and_result145[206]^and_result145[207]^and_result145[208]^and_result145[209]^and_result145[210]^and_result145[211]^and_result145[212]^and_result145[213]^and_result145[214]^and_result145[215]^and_result145[216]^and_result145[217]^and_result145[218]^and_result145[219]^and_result145[220]^and_result145[221]^and_result145[222]^and_result145[223]^and_result145[224]^and_result145[225]^and_result145[226]^and_result145[227]^and_result145[228]^and_result145[229]^and_result145[230]^and_result145[231]^and_result145[232]^and_result145[233]^and_result145[234]^and_result145[235]^and_result145[236]^and_result145[237]^and_result145[238]^and_result145[239]^and_result145[240]^and_result145[241]^and_result145[242]^and_result145[243]^and_result145[244]^and_result145[245]^and_result145[246]^and_result145[247]^and_result145[248]^and_result145[249]^and_result145[250]^and_result145[251]^and_result145[252]^and_result145[253]^and_result145[254];
assign key[146]=and_result146[0]^and_result146[1]^and_result146[2]^and_result146[3]^and_result146[4]^and_result146[5]^and_result146[6]^and_result146[7]^and_result146[8]^and_result146[9]^and_result146[10]^and_result146[11]^and_result146[12]^and_result146[13]^and_result146[14]^and_result146[15]^and_result146[16]^and_result146[17]^and_result146[18]^and_result146[19]^and_result146[20]^and_result146[21]^and_result146[22]^and_result146[23]^and_result146[24]^and_result146[25]^and_result146[26]^and_result146[27]^and_result146[28]^and_result146[29]^and_result146[30]^and_result146[31]^and_result146[32]^and_result146[33]^and_result146[34]^and_result146[35]^and_result146[36]^and_result146[37]^and_result146[38]^and_result146[39]^and_result146[40]^and_result146[41]^and_result146[42]^and_result146[43]^and_result146[44]^and_result146[45]^and_result146[46]^and_result146[47]^and_result146[48]^and_result146[49]^and_result146[50]^and_result146[51]^and_result146[52]^and_result146[53]^and_result146[54]^and_result146[55]^and_result146[56]^and_result146[57]^and_result146[58]^and_result146[59]^and_result146[60]^and_result146[61]^and_result146[62]^and_result146[63]^and_result146[64]^and_result146[65]^and_result146[66]^and_result146[67]^and_result146[68]^and_result146[69]^and_result146[70]^and_result146[71]^and_result146[72]^and_result146[73]^and_result146[74]^and_result146[75]^and_result146[76]^and_result146[77]^and_result146[78]^and_result146[79]^and_result146[80]^and_result146[81]^and_result146[82]^and_result146[83]^and_result146[84]^and_result146[85]^and_result146[86]^and_result146[87]^and_result146[88]^and_result146[89]^and_result146[90]^and_result146[91]^and_result146[92]^and_result146[93]^and_result146[94]^and_result146[95]^and_result146[96]^and_result146[97]^and_result146[98]^and_result146[99]^and_result146[100]^and_result146[101]^and_result146[102]^and_result146[103]^and_result146[104]^and_result146[105]^and_result146[106]^and_result146[107]^and_result146[108]^and_result146[109]^and_result146[110]^and_result146[111]^and_result146[112]^and_result146[113]^and_result146[114]^and_result146[115]^and_result146[116]^and_result146[117]^and_result146[118]^and_result146[119]^and_result146[120]^and_result146[121]^and_result146[122]^and_result146[123]^and_result146[124]^and_result146[125]^and_result146[126]^and_result146[127]^and_result146[128]^and_result146[129]^and_result146[130]^and_result146[131]^and_result146[132]^and_result146[133]^and_result146[134]^and_result146[135]^and_result146[136]^and_result146[137]^and_result146[138]^and_result146[139]^and_result146[140]^and_result146[141]^and_result146[142]^and_result146[143]^and_result146[144]^and_result146[145]^and_result146[146]^and_result146[147]^and_result146[148]^and_result146[149]^and_result146[150]^and_result146[151]^and_result146[152]^and_result146[153]^and_result146[154]^and_result146[155]^and_result146[156]^and_result146[157]^and_result146[158]^and_result146[159]^and_result146[160]^and_result146[161]^and_result146[162]^and_result146[163]^and_result146[164]^and_result146[165]^and_result146[166]^and_result146[167]^and_result146[168]^and_result146[169]^and_result146[170]^and_result146[171]^and_result146[172]^and_result146[173]^and_result146[174]^and_result146[175]^and_result146[176]^and_result146[177]^and_result146[178]^and_result146[179]^and_result146[180]^and_result146[181]^and_result146[182]^and_result146[183]^and_result146[184]^and_result146[185]^and_result146[186]^and_result146[187]^and_result146[188]^and_result146[189]^and_result146[190]^and_result146[191]^and_result146[192]^and_result146[193]^and_result146[194]^and_result146[195]^and_result146[196]^and_result146[197]^and_result146[198]^and_result146[199]^and_result146[200]^and_result146[201]^and_result146[202]^and_result146[203]^and_result146[204]^and_result146[205]^and_result146[206]^and_result146[207]^and_result146[208]^and_result146[209]^and_result146[210]^and_result146[211]^and_result146[212]^and_result146[213]^and_result146[214]^and_result146[215]^and_result146[216]^and_result146[217]^and_result146[218]^and_result146[219]^and_result146[220]^and_result146[221]^and_result146[222]^and_result146[223]^and_result146[224]^and_result146[225]^and_result146[226]^and_result146[227]^and_result146[228]^and_result146[229]^and_result146[230]^and_result146[231]^and_result146[232]^and_result146[233]^and_result146[234]^and_result146[235]^and_result146[236]^and_result146[237]^and_result146[238]^and_result146[239]^and_result146[240]^and_result146[241]^and_result146[242]^and_result146[243]^and_result146[244]^and_result146[245]^and_result146[246]^and_result146[247]^and_result146[248]^and_result146[249]^and_result146[250]^and_result146[251]^and_result146[252]^and_result146[253]^and_result146[254];
assign key[147]=and_result147[0]^and_result147[1]^and_result147[2]^and_result147[3]^and_result147[4]^and_result147[5]^and_result147[6]^and_result147[7]^and_result147[8]^and_result147[9]^and_result147[10]^and_result147[11]^and_result147[12]^and_result147[13]^and_result147[14]^and_result147[15]^and_result147[16]^and_result147[17]^and_result147[18]^and_result147[19]^and_result147[20]^and_result147[21]^and_result147[22]^and_result147[23]^and_result147[24]^and_result147[25]^and_result147[26]^and_result147[27]^and_result147[28]^and_result147[29]^and_result147[30]^and_result147[31]^and_result147[32]^and_result147[33]^and_result147[34]^and_result147[35]^and_result147[36]^and_result147[37]^and_result147[38]^and_result147[39]^and_result147[40]^and_result147[41]^and_result147[42]^and_result147[43]^and_result147[44]^and_result147[45]^and_result147[46]^and_result147[47]^and_result147[48]^and_result147[49]^and_result147[50]^and_result147[51]^and_result147[52]^and_result147[53]^and_result147[54]^and_result147[55]^and_result147[56]^and_result147[57]^and_result147[58]^and_result147[59]^and_result147[60]^and_result147[61]^and_result147[62]^and_result147[63]^and_result147[64]^and_result147[65]^and_result147[66]^and_result147[67]^and_result147[68]^and_result147[69]^and_result147[70]^and_result147[71]^and_result147[72]^and_result147[73]^and_result147[74]^and_result147[75]^and_result147[76]^and_result147[77]^and_result147[78]^and_result147[79]^and_result147[80]^and_result147[81]^and_result147[82]^and_result147[83]^and_result147[84]^and_result147[85]^and_result147[86]^and_result147[87]^and_result147[88]^and_result147[89]^and_result147[90]^and_result147[91]^and_result147[92]^and_result147[93]^and_result147[94]^and_result147[95]^and_result147[96]^and_result147[97]^and_result147[98]^and_result147[99]^and_result147[100]^and_result147[101]^and_result147[102]^and_result147[103]^and_result147[104]^and_result147[105]^and_result147[106]^and_result147[107]^and_result147[108]^and_result147[109]^and_result147[110]^and_result147[111]^and_result147[112]^and_result147[113]^and_result147[114]^and_result147[115]^and_result147[116]^and_result147[117]^and_result147[118]^and_result147[119]^and_result147[120]^and_result147[121]^and_result147[122]^and_result147[123]^and_result147[124]^and_result147[125]^and_result147[126]^and_result147[127]^and_result147[128]^and_result147[129]^and_result147[130]^and_result147[131]^and_result147[132]^and_result147[133]^and_result147[134]^and_result147[135]^and_result147[136]^and_result147[137]^and_result147[138]^and_result147[139]^and_result147[140]^and_result147[141]^and_result147[142]^and_result147[143]^and_result147[144]^and_result147[145]^and_result147[146]^and_result147[147]^and_result147[148]^and_result147[149]^and_result147[150]^and_result147[151]^and_result147[152]^and_result147[153]^and_result147[154]^and_result147[155]^and_result147[156]^and_result147[157]^and_result147[158]^and_result147[159]^and_result147[160]^and_result147[161]^and_result147[162]^and_result147[163]^and_result147[164]^and_result147[165]^and_result147[166]^and_result147[167]^and_result147[168]^and_result147[169]^and_result147[170]^and_result147[171]^and_result147[172]^and_result147[173]^and_result147[174]^and_result147[175]^and_result147[176]^and_result147[177]^and_result147[178]^and_result147[179]^and_result147[180]^and_result147[181]^and_result147[182]^and_result147[183]^and_result147[184]^and_result147[185]^and_result147[186]^and_result147[187]^and_result147[188]^and_result147[189]^and_result147[190]^and_result147[191]^and_result147[192]^and_result147[193]^and_result147[194]^and_result147[195]^and_result147[196]^and_result147[197]^and_result147[198]^and_result147[199]^and_result147[200]^and_result147[201]^and_result147[202]^and_result147[203]^and_result147[204]^and_result147[205]^and_result147[206]^and_result147[207]^and_result147[208]^and_result147[209]^and_result147[210]^and_result147[211]^and_result147[212]^and_result147[213]^and_result147[214]^and_result147[215]^and_result147[216]^and_result147[217]^and_result147[218]^and_result147[219]^and_result147[220]^and_result147[221]^and_result147[222]^and_result147[223]^and_result147[224]^and_result147[225]^and_result147[226]^and_result147[227]^and_result147[228]^and_result147[229]^and_result147[230]^and_result147[231]^and_result147[232]^and_result147[233]^and_result147[234]^and_result147[235]^and_result147[236]^and_result147[237]^and_result147[238]^and_result147[239]^and_result147[240]^and_result147[241]^and_result147[242]^and_result147[243]^and_result147[244]^and_result147[245]^and_result147[246]^and_result147[247]^and_result147[248]^and_result147[249]^and_result147[250]^and_result147[251]^and_result147[252]^and_result147[253]^and_result147[254];
assign key[148]=and_result148[0]^and_result148[1]^and_result148[2]^and_result148[3]^and_result148[4]^and_result148[5]^and_result148[6]^and_result148[7]^and_result148[8]^and_result148[9]^and_result148[10]^and_result148[11]^and_result148[12]^and_result148[13]^and_result148[14]^and_result148[15]^and_result148[16]^and_result148[17]^and_result148[18]^and_result148[19]^and_result148[20]^and_result148[21]^and_result148[22]^and_result148[23]^and_result148[24]^and_result148[25]^and_result148[26]^and_result148[27]^and_result148[28]^and_result148[29]^and_result148[30]^and_result148[31]^and_result148[32]^and_result148[33]^and_result148[34]^and_result148[35]^and_result148[36]^and_result148[37]^and_result148[38]^and_result148[39]^and_result148[40]^and_result148[41]^and_result148[42]^and_result148[43]^and_result148[44]^and_result148[45]^and_result148[46]^and_result148[47]^and_result148[48]^and_result148[49]^and_result148[50]^and_result148[51]^and_result148[52]^and_result148[53]^and_result148[54]^and_result148[55]^and_result148[56]^and_result148[57]^and_result148[58]^and_result148[59]^and_result148[60]^and_result148[61]^and_result148[62]^and_result148[63]^and_result148[64]^and_result148[65]^and_result148[66]^and_result148[67]^and_result148[68]^and_result148[69]^and_result148[70]^and_result148[71]^and_result148[72]^and_result148[73]^and_result148[74]^and_result148[75]^and_result148[76]^and_result148[77]^and_result148[78]^and_result148[79]^and_result148[80]^and_result148[81]^and_result148[82]^and_result148[83]^and_result148[84]^and_result148[85]^and_result148[86]^and_result148[87]^and_result148[88]^and_result148[89]^and_result148[90]^and_result148[91]^and_result148[92]^and_result148[93]^and_result148[94]^and_result148[95]^and_result148[96]^and_result148[97]^and_result148[98]^and_result148[99]^and_result148[100]^and_result148[101]^and_result148[102]^and_result148[103]^and_result148[104]^and_result148[105]^and_result148[106]^and_result148[107]^and_result148[108]^and_result148[109]^and_result148[110]^and_result148[111]^and_result148[112]^and_result148[113]^and_result148[114]^and_result148[115]^and_result148[116]^and_result148[117]^and_result148[118]^and_result148[119]^and_result148[120]^and_result148[121]^and_result148[122]^and_result148[123]^and_result148[124]^and_result148[125]^and_result148[126]^and_result148[127]^and_result148[128]^and_result148[129]^and_result148[130]^and_result148[131]^and_result148[132]^and_result148[133]^and_result148[134]^and_result148[135]^and_result148[136]^and_result148[137]^and_result148[138]^and_result148[139]^and_result148[140]^and_result148[141]^and_result148[142]^and_result148[143]^and_result148[144]^and_result148[145]^and_result148[146]^and_result148[147]^and_result148[148]^and_result148[149]^and_result148[150]^and_result148[151]^and_result148[152]^and_result148[153]^and_result148[154]^and_result148[155]^and_result148[156]^and_result148[157]^and_result148[158]^and_result148[159]^and_result148[160]^and_result148[161]^and_result148[162]^and_result148[163]^and_result148[164]^and_result148[165]^and_result148[166]^and_result148[167]^and_result148[168]^and_result148[169]^and_result148[170]^and_result148[171]^and_result148[172]^and_result148[173]^and_result148[174]^and_result148[175]^and_result148[176]^and_result148[177]^and_result148[178]^and_result148[179]^and_result148[180]^and_result148[181]^and_result148[182]^and_result148[183]^and_result148[184]^and_result148[185]^and_result148[186]^and_result148[187]^and_result148[188]^and_result148[189]^and_result148[190]^and_result148[191]^and_result148[192]^and_result148[193]^and_result148[194]^and_result148[195]^and_result148[196]^and_result148[197]^and_result148[198]^and_result148[199]^and_result148[200]^and_result148[201]^and_result148[202]^and_result148[203]^and_result148[204]^and_result148[205]^and_result148[206]^and_result148[207]^and_result148[208]^and_result148[209]^and_result148[210]^and_result148[211]^and_result148[212]^and_result148[213]^and_result148[214]^and_result148[215]^and_result148[216]^and_result148[217]^and_result148[218]^and_result148[219]^and_result148[220]^and_result148[221]^and_result148[222]^and_result148[223]^and_result148[224]^and_result148[225]^and_result148[226]^and_result148[227]^and_result148[228]^and_result148[229]^and_result148[230]^and_result148[231]^and_result148[232]^and_result148[233]^and_result148[234]^and_result148[235]^and_result148[236]^and_result148[237]^and_result148[238]^and_result148[239]^and_result148[240]^and_result148[241]^and_result148[242]^and_result148[243]^and_result148[244]^and_result148[245]^and_result148[246]^and_result148[247]^and_result148[248]^and_result148[249]^and_result148[250]^and_result148[251]^and_result148[252]^and_result148[253]^and_result148[254];
assign key[149]=and_result149[0]^and_result149[1]^and_result149[2]^and_result149[3]^and_result149[4]^and_result149[5]^and_result149[6]^and_result149[7]^and_result149[8]^and_result149[9]^and_result149[10]^and_result149[11]^and_result149[12]^and_result149[13]^and_result149[14]^and_result149[15]^and_result149[16]^and_result149[17]^and_result149[18]^and_result149[19]^and_result149[20]^and_result149[21]^and_result149[22]^and_result149[23]^and_result149[24]^and_result149[25]^and_result149[26]^and_result149[27]^and_result149[28]^and_result149[29]^and_result149[30]^and_result149[31]^and_result149[32]^and_result149[33]^and_result149[34]^and_result149[35]^and_result149[36]^and_result149[37]^and_result149[38]^and_result149[39]^and_result149[40]^and_result149[41]^and_result149[42]^and_result149[43]^and_result149[44]^and_result149[45]^and_result149[46]^and_result149[47]^and_result149[48]^and_result149[49]^and_result149[50]^and_result149[51]^and_result149[52]^and_result149[53]^and_result149[54]^and_result149[55]^and_result149[56]^and_result149[57]^and_result149[58]^and_result149[59]^and_result149[60]^and_result149[61]^and_result149[62]^and_result149[63]^and_result149[64]^and_result149[65]^and_result149[66]^and_result149[67]^and_result149[68]^and_result149[69]^and_result149[70]^and_result149[71]^and_result149[72]^and_result149[73]^and_result149[74]^and_result149[75]^and_result149[76]^and_result149[77]^and_result149[78]^and_result149[79]^and_result149[80]^and_result149[81]^and_result149[82]^and_result149[83]^and_result149[84]^and_result149[85]^and_result149[86]^and_result149[87]^and_result149[88]^and_result149[89]^and_result149[90]^and_result149[91]^and_result149[92]^and_result149[93]^and_result149[94]^and_result149[95]^and_result149[96]^and_result149[97]^and_result149[98]^and_result149[99]^and_result149[100]^and_result149[101]^and_result149[102]^and_result149[103]^and_result149[104]^and_result149[105]^and_result149[106]^and_result149[107]^and_result149[108]^and_result149[109]^and_result149[110]^and_result149[111]^and_result149[112]^and_result149[113]^and_result149[114]^and_result149[115]^and_result149[116]^and_result149[117]^and_result149[118]^and_result149[119]^and_result149[120]^and_result149[121]^and_result149[122]^and_result149[123]^and_result149[124]^and_result149[125]^and_result149[126]^and_result149[127]^and_result149[128]^and_result149[129]^and_result149[130]^and_result149[131]^and_result149[132]^and_result149[133]^and_result149[134]^and_result149[135]^and_result149[136]^and_result149[137]^and_result149[138]^and_result149[139]^and_result149[140]^and_result149[141]^and_result149[142]^and_result149[143]^and_result149[144]^and_result149[145]^and_result149[146]^and_result149[147]^and_result149[148]^and_result149[149]^and_result149[150]^and_result149[151]^and_result149[152]^and_result149[153]^and_result149[154]^and_result149[155]^and_result149[156]^and_result149[157]^and_result149[158]^and_result149[159]^and_result149[160]^and_result149[161]^and_result149[162]^and_result149[163]^and_result149[164]^and_result149[165]^and_result149[166]^and_result149[167]^and_result149[168]^and_result149[169]^and_result149[170]^and_result149[171]^and_result149[172]^and_result149[173]^and_result149[174]^and_result149[175]^and_result149[176]^and_result149[177]^and_result149[178]^and_result149[179]^and_result149[180]^and_result149[181]^and_result149[182]^and_result149[183]^and_result149[184]^and_result149[185]^and_result149[186]^and_result149[187]^and_result149[188]^and_result149[189]^and_result149[190]^and_result149[191]^and_result149[192]^and_result149[193]^and_result149[194]^and_result149[195]^and_result149[196]^and_result149[197]^and_result149[198]^and_result149[199]^and_result149[200]^and_result149[201]^and_result149[202]^and_result149[203]^and_result149[204]^and_result149[205]^and_result149[206]^and_result149[207]^and_result149[208]^and_result149[209]^and_result149[210]^and_result149[211]^and_result149[212]^and_result149[213]^and_result149[214]^and_result149[215]^and_result149[216]^and_result149[217]^and_result149[218]^and_result149[219]^and_result149[220]^and_result149[221]^and_result149[222]^and_result149[223]^and_result149[224]^and_result149[225]^and_result149[226]^and_result149[227]^and_result149[228]^and_result149[229]^and_result149[230]^and_result149[231]^and_result149[232]^and_result149[233]^and_result149[234]^and_result149[235]^and_result149[236]^and_result149[237]^and_result149[238]^and_result149[239]^and_result149[240]^and_result149[241]^and_result149[242]^and_result149[243]^and_result149[244]^and_result149[245]^and_result149[246]^and_result149[247]^and_result149[248]^and_result149[249]^and_result149[250]^and_result149[251]^and_result149[252]^and_result149[253]^and_result149[254];
assign key[150]=and_result150[0]^and_result150[1]^and_result150[2]^and_result150[3]^and_result150[4]^and_result150[5]^and_result150[6]^and_result150[7]^and_result150[8]^and_result150[9]^and_result150[10]^and_result150[11]^and_result150[12]^and_result150[13]^and_result150[14]^and_result150[15]^and_result150[16]^and_result150[17]^and_result150[18]^and_result150[19]^and_result150[20]^and_result150[21]^and_result150[22]^and_result150[23]^and_result150[24]^and_result150[25]^and_result150[26]^and_result150[27]^and_result150[28]^and_result150[29]^and_result150[30]^and_result150[31]^and_result150[32]^and_result150[33]^and_result150[34]^and_result150[35]^and_result150[36]^and_result150[37]^and_result150[38]^and_result150[39]^and_result150[40]^and_result150[41]^and_result150[42]^and_result150[43]^and_result150[44]^and_result150[45]^and_result150[46]^and_result150[47]^and_result150[48]^and_result150[49]^and_result150[50]^and_result150[51]^and_result150[52]^and_result150[53]^and_result150[54]^and_result150[55]^and_result150[56]^and_result150[57]^and_result150[58]^and_result150[59]^and_result150[60]^and_result150[61]^and_result150[62]^and_result150[63]^and_result150[64]^and_result150[65]^and_result150[66]^and_result150[67]^and_result150[68]^and_result150[69]^and_result150[70]^and_result150[71]^and_result150[72]^and_result150[73]^and_result150[74]^and_result150[75]^and_result150[76]^and_result150[77]^and_result150[78]^and_result150[79]^and_result150[80]^and_result150[81]^and_result150[82]^and_result150[83]^and_result150[84]^and_result150[85]^and_result150[86]^and_result150[87]^and_result150[88]^and_result150[89]^and_result150[90]^and_result150[91]^and_result150[92]^and_result150[93]^and_result150[94]^and_result150[95]^and_result150[96]^and_result150[97]^and_result150[98]^and_result150[99]^and_result150[100]^and_result150[101]^and_result150[102]^and_result150[103]^and_result150[104]^and_result150[105]^and_result150[106]^and_result150[107]^and_result150[108]^and_result150[109]^and_result150[110]^and_result150[111]^and_result150[112]^and_result150[113]^and_result150[114]^and_result150[115]^and_result150[116]^and_result150[117]^and_result150[118]^and_result150[119]^and_result150[120]^and_result150[121]^and_result150[122]^and_result150[123]^and_result150[124]^and_result150[125]^and_result150[126]^and_result150[127]^and_result150[128]^and_result150[129]^and_result150[130]^and_result150[131]^and_result150[132]^and_result150[133]^and_result150[134]^and_result150[135]^and_result150[136]^and_result150[137]^and_result150[138]^and_result150[139]^and_result150[140]^and_result150[141]^and_result150[142]^and_result150[143]^and_result150[144]^and_result150[145]^and_result150[146]^and_result150[147]^and_result150[148]^and_result150[149]^and_result150[150]^and_result150[151]^and_result150[152]^and_result150[153]^and_result150[154]^and_result150[155]^and_result150[156]^and_result150[157]^and_result150[158]^and_result150[159]^and_result150[160]^and_result150[161]^and_result150[162]^and_result150[163]^and_result150[164]^and_result150[165]^and_result150[166]^and_result150[167]^and_result150[168]^and_result150[169]^and_result150[170]^and_result150[171]^and_result150[172]^and_result150[173]^and_result150[174]^and_result150[175]^and_result150[176]^and_result150[177]^and_result150[178]^and_result150[179]^and_result150[180]^and_result150[181]^and_result150[182]^and_result150[183]^and_result150[184]^and_result150[185]^and_result150[186]^and_result150[187]^and_result150[188]^and_result150[189]^and_result150[190]^and_result150[191]^and_result150[192]^and_result150[193]^and_result150[194]^and_result150[195]^and_result150[196]^and_result150[197]^and_result150[198]^and_result150[199]^and_result150[200]^and_result150[201]^and_result150[202]^and_result150[203]^and_result150[204]^and_result150[205]^and_result150[206]^and_result150[207]^and_result150[208]^and_result150[209]^and_result150[210]^and_result150[211]^and_result150[212]^and_result150[213]^and_result150[214]^and_result150[215]^and_result150[216]^and_result150[217]^and_result150[218]^and_result150[219]^and_result150[220]^and_result150[221]^and_result150[222]^and_result150[223]^and_result150[224]^and_result150[225]^and_result150[226]^and_result150[227]^and_result150[228]^and_result150[229]^and_result150[230]^and_result150[231]^and_result150[232]^and_result150[233]^and_result150[234]^and_result150[235]^and_result150[236]^and_result150[237]^and_result150[238]^and_result150[239]^and_result150[240]^and_result150[241]^and_result150[242]^and_result150[243]^and_result150[244]^and_result150[245]^and_result150[246]^and_result150[247]^and_result150[248]^and_result150[249]^and_result150[250]^and_result150[251]^and_result150[252]^and_result150[253]^and_result150[254];
assign key[151]=and_result151[0]^and_result151[1]^and_result151[2]^and_result151[3]^and_result151[4]^and_result151[5]^and_result151[6]^and_result151[7]^and_result151[8]^and_result151[9]^and_result151[10]^and_result151[11]^and_result151[12]^and_result151[13]^and_result151[14]^and_result151[15]^and_result151[16]^and_result151[17]^and_result151[18]^and_result151[19]^and_result151[20]^and_result151[21]^and_result151[22]^and_result151[23]^and_result151[24]^and_result151[25]^and_result151[26]^and_result151[27]^and_result151[28]^and_result151[29]^and_result151[30]^and_result151[31]^and_result151[32]^and_result151[33]^and_result151[34]^and_result151[35]^and_result151[36]^and_result151[37]^and_result151[38]^and_result151[39]^and_result151[40]^and_result151[41]^and_result151[42]^and_result151[43]^and_result151[44]^and_result151[45]^and_result151[46]^and_result151[47]^and_result151[48]^and_result151[49]^and_result151[50]^and_result151[51]^and_result151[52]^and_result151[53]^and_result151[54]^and_result151[55]^and_result151[56]^and_result151[57]^and_result151[58]^and_result151[59]^and_result151[60]^and_result151[61]^and_result151[62]^and_result151[63]^and_result151[64]^and_result151[65]^and_result151[66]^and_result151[67]^and_result151[68]^and_result151[69]^and_result151[70]^and_result151[71]^and_result151[72]^and_result151[73]^and_result151[74]^and_result151[75]^and_result151[76]^and_result151[77]^and_result151[78]^and_result151[79]^and_result151[80]^and_result151[81]^and_result151[82]^and_result151[83]^and_result151[84]^and_result151[85]^and_result151[86]^and_result151[87]^and_result151[88]^and_result151[89]^and_result151[90]^and_result151[91]^and_result151[92]^and_result151[93]^and_result151[94]^and_result151[95]^and_result151[96]^and_result151[97]^and_result151[98]^and_result151[99]^and_result151[100]^and_result151[101]^and_result151[102]^and_result151[103]^and_result151[104]^and_result151[105]^and_result151[106]^and_result151[107]^and_result151[108]^and_result151[109]^and_result151[110]^and_result151[111]^and_result151[112]^and_result151[113]^and_result151[114]^and_result151[115]^and_result151[116]^and_result151[117]^and_result151[118]^and_result151[119]^and_result151[120]^and_result151[121]^and_result151[122]^and_result151[123]^and_result151[124]^and_result151[125]^and_result151[126]^and_result151[127]^and_result151[128]^and_result151[129]^and_result151[130]^and_result151[131]^and_result151[132]^and_result151[133]^and_result151[134]^and_result151[135]^and_result151[136]^and_result151[137]^and_result151[138]^and_result151[139]^and_result151[140]^and_result151[141]^and_result151[142]^and_result151[143]^and_result151[144]^and_result151[145]^and_result151[146]^and_result151[147]^and_result151[148]^and_result151[149]^and_result151[150]^and_result151[151]^and_result151[152]^and_result151[153]^and_result151[154]^and_result151[155]^and_result151[156]^and_result151[157]^and_result151[158]^and_result151[159]^and_result151[160]^and_result151[161]^and_result151[162]^and_result151[163]^and_result151[164]^and_result151[165]^and_result151[166]^and_result151[167]^and_result151[168]^and_result151[169]^and_result151[170]^and_result151[171]^and_result151[172]^and_result151[173]^and_result151[174]^and_result151[175]^and_result151[176]^and_result151[177]^and_result151[178]^and_result151[179]^and_result151[180]^and_result151[181]^and_result151[182]^and_result151[183]^and_result151[184]^and_result151[185]^and_result151[186]^and_result151[187]^and_result151[188]^and_result151[189]^and_result151[190]^and_result151[191]^and_result151[192]^and_result151[193]^and_result151[194]^and_result151[195]^and_result151[196]^and_result151[197]^and_result151[198]^and_result151[199]^and_result151[200]^and_result151[201]^and_result151[202]^and_result151[203]^and_result151[204]^and_result151[205]^and_result151[206]^and_result151[207]^and_result151[208]^and_result151[209]^and_result151[210]^and_result151[211]^and_result151[212]^and_result151[213]^and_result151[214]^and_result151[215]^and_result151[216]^and_result151[217]^and_result151[218]^and_result151[219]^and_result151[220]^and_result151[221]^and_result151[222]^and_result151[223]^and_result151[224]^and_result151[225]^and_result151[226]^and_result151[227]^and_result151[228]^and_result151[229]^and_result151[230]^and_result151[231]^and_result151[232]^and_result151[233]^and_result151[234]^and_result151[235]^and_result151[236]^and_result151[237]^and_result151[238]^and_result151[239]^and_result151[240]^and_result151[241]^and_result151[242]^and_result151[243]^and_result151[244]^and_result151[245]^and_result151[246]^and_result151[247]^and_result151[248]^and_result151[249]^and_result151[250]^and_result151[251]^and_result151[252]^and_result151[253]^and_result151[254];
assign key[152]=and_result152[0]^and_result152[1]^and_result152[2]^and_result152[3]^and_result152[4]^and_result152[5]^and_result152[6]^and_result152[7]^and_result152[8]^and_result152[9]^and_result152[10]^and_result152[11]^and_result152[12]^and_result152[13]^and_result152[14]^and_result152[15]^and_result152[16]^and_result152[17]^and_result152[18]^and_result152[19]^and_result152[20]^and_result152[21]^and_result152[22]^and_result152[23]^and_result152[24]^and_result152[25]^and_result152[26]^and_result152[27]^and_result152[28]^and_result152[29]^and_result152[30]^and_result152[31]^and_result152[32]^and_result152[33]^and_result152[34]^and_result152[35]^and_result152[36]^and_result152[37]^and_result152[38]^and_result152[39]^and_result152[40]^and_result152[41]^and_result152[42]^and_result152[43]^and_result152[44]^and_result152[45]^and_result152[46]^and_result152[47]^and_result152[48]^and_result152[49]^and_result152[50]^and_result152[51]^and_result152[52]^and_result152[53]^and_result152[54]^and_result152[55]^and_result152[56]^and_result152[57]^and_result152[58]^and_result152[59]^and_result152[60]^and_result152[61]^and_result152[62]^and_result152[63]^and_result152[64]^and_result152[65]^and_result152[66]^and_result152[67]^and_result152[68]^and_result152[69]^and_result152[70]^and_result152[71]^and_result152[72]^and_result152[73]^and_result152[74]^and_result152[75]^and_result152[76]^and_result152[77]^and_result152[78]^and_result152[79]^and_result152[80]^and_result152[81]^and_result152[82]^and_result152[83]^and_result152[84]^and_result152[85]^and_result152[86]^and_result152[87]^and_result152[88]^and_result152[89]^and_result152[90]^and_result152[91]^and_result152[92]^and_result152[93]^and_result152[94]^and_result152[95]^and_result152[96]^and_result152[97]^and_result152[98]^and_result152[99]^and_result152[100]^and_result152[101]^and_result152[102]^and_result152[103]^and_result152[104]^and_result152[105]^and_result152[106]^and_result152[107]^and_result152[108]^and_result152[109]^and_result152[110]^and_result152[111]^and_result152[112]^and_result152[113]^and_result152[114]^and_result152[115]^and_result152[116]^and_result152[117]^and_result152[118]^and_result152[119]^and_result152[120]^and_result152[121]^and_result152[122]^and_result152[123]^and_result152[124]^and_result152[125]^and_result152[126]^and_result152[127]^and_result152[128]^and_result152[129]^and_result152[130]^and_result152[131]^and_result152[132]^and_result152[133]^and_result152[134]^and_result152[135]^and_result152[136]^and_result152[137]^and_result152[138]^and_result152[139]^and_result152[140]^and_result152[141]^and_result152[142]^and_result152[143]^and_result152[144]^and_result152[145]^and_result152[146]^and_result152[147]^and_result152[148]^and_result152[149]^and_result152[150]^and_result152[151]^and_result152[152]^and_result152[153]^and_result152[154]^and_result152[155]^and_result152[156]^and_result152[157]^and_result152[158]^and_result152[159]^and_result152[160]^and_result152[161]^and_result152[162]^and_result152[163]^and_result152[164]^and_result152[165]^and_result152[166]^and_result152[167]^and_result152[168]^and_result152[169]^and_result152[170]^and_result152[171]^and_result152[172]^and_result152[173]^and_result152[174]^and_result152[175]^and_result152[176]^and_result152[177]^and_result152[178]^and_result152[179]^and_result152[180]^and_result152[181]^and_result152[182]^and_result152[183]^and_result152[184]^and_result152[185]^and_result152[186]^and_result152[187]^and_result152[188]^and_result152[189]^and_result152[190]^and_result152[191]^and_result152[192]^and_result152[193]^and_result152[194]^and_result152[195]^and_result152[196]^and_result152[197]^and_result152[198]^and_result152[199]^and_result152[200]^and_result152[201]^and_result152[202]^and_result152[203]^and_result152[204]^and_result152[205]^and_result152[206]^and_result152[207]^and_result152[208]^and_result152[209]^and_result152[210]^and_result152[211]^and_result152[212]^and_result152[213]^and_result152[214]^and_result152[215]^and_result152[216]^and_result152[217]^and_result152[218]^and_result152[219]^and_result152[220]^and_result152[221]^and_result152[222]^and_result152[223]^and_result152[224]^and_result152[225]^and_result152[226]^and_result152[227]^and_result152[228]^and_result152[229]^and_result152[230]^and_result152[231]^and_result152[232]^and_result152[233]^and_result152[234]^and_result152[235]^and_result152[236]^and_result152[237]^and_result152[238]^and_result152[239]^and_result152[240]^and_result152[241]^and_result152[242]^and_result152[243]^and_result152[244]^and_result152[245]^and_result152[246]^and_result152[247]^and_result152[248]^and_result152[249]^and_result152[250]^and_result152[251]^and_result152[252]^and_result152[253]^and_result152[254];
assign key[153]=and_result153[0]^and_result153[1]^and_result153[2]^and_result153[3]^and_result153[4]^and_result153[5]^and_result153[6]^and_result153[7]^and_result153[8]^and_result153[9]^and_result153[10]^and_result153[11]^and_result153[12]^and_result153[13]^and_result153[14]^and_result153[15]^and_result153[16]^and_result153[17]^and_result153[18]^and_result153[19]^and_result153[20]^and_result153[21]^and_result153[22]^and_result153[23]^and_result153[24]^and_result153[25]^and_result153[26]^and_result153[27]^and_result153[28]^and_result153[29]^and_result153[30]^and_result153[31]^and_result153[32]^and_result153[33]^and_result153[34]^and_result153[35]^and_result153[36]^and_result153[37]^and_result153[38]^and_result153[39]^and_result153[40]^and_result153[41]^and_result153[42]^and_result153[43]^and_result153[44]^and_result153[45]^and_result153[46]^and_result153[47]^and_result153[48]^and_result153[49]^and_result153[50]^and_result153[51]^and_result153[52]^and_result153[53]^and_result153[54]^and_result153[55]^and_result153[56]^and_result153[57]^and_result153[58]^and_result153[59]^and_result153[60]^and_result153[61]^and_result153[62]^and_result153[63]^and_result153[64]^and_result153[65]^and_result153[66]^and_result153[67]^and_result153[68]^and_result153[69]^and_result153[70]^and_result153[71]^and_result153[72]^and_result153[73]^and_result153[74]^and_result153[75]^and_result153[76]^and_result153[77]^and_result153[78]^and_result153[79]^and_result153[80]^and_result153[81]^and_result153[82]^and_result153[83]^and_result153[84]^and_result153[85]^and_result153[86]^and_result153[87]^and_result153[88]^and_result153[89]^and_result153[90]^and_result153[91]^and_result153[92]^and_result153[93]^and_result153[94]^and_result153[95]^and_result153[96]^and_result153[97]^and_result153[98]^and_result153[99]^and_result153[100]^and_result153[101]^and_result153[102]^and_result153[103]^and_result153[104]^and_result153[105]^and_result153[106]^and_result153[107]^and_result153[108]^and_result153[109]^and_result153[110]^and_result153[111]^and_result153[112]^and_result153[113]^and_result153[114]^and_result153[115]^and_result153[116]^and_result153[117]^and_result153[118]^and_result153[119]^and_result153[120]^and_result153[121]^and_result153[122]^and_result153[123]^and_result153[124]^and_result153[125]^and_result153[126]^and_result153[127]^and_result153[128]^and_result153[129]^and_result153[130]^and_result153[131]^and_result153[132]^and_result153[133]^and_result153[134]^and_result153[135]^and_result153[136]^and_result153[137]^and_result153[138]^and_result153[139]^and_result153[140]^and_result153[141]^and_result153[142]^and_result153[143]^and_result153[144]^and_result153[145]^and_result153[146]^and_result153[147]^and_result153[148]^and_result153[149]^and_result153[150]^and_result153[151]^and_result153[152]^and_result153[153]^and_result153[154]^and_result153[155]^and_result153[156]^and_result153[157]^and_result153[158]^and_result153[159]^and_result153[160]^and_result153[161]^and_result153[162]^and_result153[163]^and_result153[164]^and_result153[165]^and_result153[166]^and_result153[167]^and_result153[168]^and_result153[169]^and_result153[170]^and_result153[171]^and_result153[172]^and_result153[173]^and_result153[174]^and_result153[175]^and_result153[176]^and_result153[177]^and_result153[178]^and_result153[179]^and_result153[180]^and_result153[181]^and_result153[182]^and_result153[183]^and_result153[184]^and_result153[185]^and_result153[186]^and_result153[187]^and_result153[188]^and_result153[189]^and_result153[190]^and_result153[191]^and_result153[192]^and_result153[193]^and_result153[194]^and_result153[195]^and_result153[196]^and_result153[197]^and_result153[198]^and_result153[199]^and_result153[200]^and_result153[201]^and_result153[202]^and_result153[203]^and_result153[204]^and_result153[205]^and_result153[206]^and_result153[207]^and_result153[208]^and_result153[209]^and_result153[210]^and_result153[211]^and_result153[212]^and_result153[213]^and_result153[214]^and_result153[215]^and_result153[216]^and_result153[217]^and_result153[218]^and_result153[219]^and_result153[220]^and_result153[221]^and_result153[222]^and_result153[223]^and_result153[224]^and_result153[225]^and_result153[226]^and_result153[227]^and_result153[228]^and_result153[229]^and_result153[230]^and_result153[231]^and_result153[232]^and_result153[233]^and_result153[234]^and_result153[235]^and_result153[236]^and_result153[237]^and_result153[238]^and_result153[239]^and_result153[240]^and_result153[241]^and_result153[242]^and_result153[243]^and_result153[244]^and_result153[245]^and_result153[246]^and_result153[247]^and_result153[248]^and_result153[249]^and_result153[250]^and_result153[251]^and_result153[252]^and_result153[253]^and_result153[254];
assign key[154]=and_result154[0]^and_result154[1]^and_result154[2]^and_result154[3]^and_result154[4]^and_result154[5]^and_result154[6]^and_result154[7]^and_result154[8]^and_result154[9]^and_result154[10]^and_result154[11]^and_result154[12]^and_result154[13]^and_result154[14]^and_result154[15]^and_result154[16]^and_result154[17]^and_result154[18]^and_result154[19]^and_result154[20]^and_result154[21]^and_result154[22]^and_result154[23]^and_result154[24]^and_result154[25]^and_result154[26]^and_result154[27]^and_result154[28]^and_result154[29]^and_result154[30]^and_result154[31]^and_result154[32]^and_result154[33]^and_result154[34]^and_result154[35]^and_result154[36]^and_result154[37]^and_result154[38]^and_result154[39]^and_result154[40]^and_result154[41]^and_result154[42]^and_result154[43]^and_result154[44]^and_result154[45]^and_result154[46]^and_result154[47]^and_result154[48]^and_result154[49]^and_result154[50]^and_result154[51]^and_result154[52]^and_result154[53]^and_result154[54]^and_result154[55]^and_result154[56]^and_result154[57]^and_result154[58]^and_result154[59]^and_result154[60]^and_result154[61]^and_result154[62]^and_result154[63]^and_result154[64]^and_result154[65]^and_result154[66]^and_result154[67]^and_result154[68]^and_result154[69]^and_result154[70]^and_result154[71]^and_result154[72]^and_result154[73]^and_result154[74]^and_result154[75]^and_result154[76]^and_result154[77]^and_result154[78]^and_result154[79]^and_result154[80]^and_result154[81]^and_result154[82]^and_result154[83]^and_result154[84]^and_result154[85]^and_result154[86]^and_result154[87]^and_result154[88]^and_result154[89]^and_result154[90]^and_result154[91]^and_result154[92]^and_result154[93]^and_result154[94]^and_result154[95]^and_result154[96]^and_result154[97]^and_result154[98]^and_result154[99]^and_result154[100]^and_result154[101]^and_result154[102]^and_result154[103]^and_result154[104]^and_result154[105]^and_result154[106]^and_result154[107]^and_result154[108]^and_result154[109]^and_result154[110]^and_result154[111]^and_result154[112]^and_result154[113]^and_result154[114]^and_result154[115]^and_result154[116]^and_result154[117]^and_result154[118]^and_result154[119]^and_result154[120]^and_result154[121]^and_result154[122]^and_result154[123]^and_result154[124]^and_result154[125]^and_result154[126]^and_result154[127]^and_result154[128]^and_result154[129]^and_result154[130]^and_result154[131]^and_result154[132]^and_result154[133]^and_result154[134]^and_result154[135]^and_result154[136]^and_result154[137]^and_result154[138]^and_result154[139]^and_result154[140]^and_result154[141]^and_result154[142]^and_result154[143]^and_result154[144]^and_result154[145]^and_result154[146]^and_result154[147]^and_result154[148]^and_result154[149]^and_result154[150]^and_result154[151]^and_result154[152]^and_result154[153]^and_result154[154]^and_result154[155]^and_result154[156]^and_result154[157]^and_result154[158]^and_result154[159]^and_result154[160]^and_result154[161]^and_result154[162]^and_result154[163]^and_result154[164]^and_result154[165]^and_result154[166]^and_result154[167]^and_result154[168]^and_result154[169]^and_result154[170]^and_result154[171]^and_result154[172]^and_result154[173]^and_result154[174]^and_result154[175]^and_result154[176]^and_result154[177]^and_result154[178]^and_result154[179]^and_result154[180]^and_result154[181]^and_result154[182]^and_result154[183]^and_result154[184]^and_result154[185]^and_result154[186]^and_result154[187]^and_result154[188]^and_result154[189]^and_result154[190]^and_result154[191]^and_result154[192]^and_result154[193]^and_result154[194]^and_result154[195]^and_result154[196]^and_result154[197]^and_result154[198]^and_result154[199]^and_result154[200]^and_result154[201]^and_result154[202]^and_result154[203]^and_result154[204]^and_result154[205]^and_result154[206]^and_result154[207]^and_result154[208]^and_result154[209]^and_result154[210]^and_result154[211]^and_result154[212]^and_result154[213]^and_result154[214]^and_result154[215]^and_result154[216]^and_result154[217]^and_result154[218]^and_result154[219]^and_result154[220]^and_result154[221]^and_result154[222]^and_result154[223]^and_result154[224]^and_result154[225]^and_result154[226]^and_result154[227]^and_result154[228]^and_result154[229]^and_result154[230]^and_result154[231]^and_result154[232]^and_result154[233]^and_result154[234]^and_result154[235]^and_result154[236]^and_result154[237]^and_result154[238]^and_result154[239]^and_result154[240]^and_result154[241]^and_result154[242]^and_result154[243]^and_result154[244]^and_result154[245]^and_result154[246]^and_result154[247]^and_result154[248]^and_result154[249]^and_result154[250]^and_result154[251]^and_result154[252]^and_result154[253]^and_result154[254];
assign key[155]=and_result155[0]^and_result155[1]^and_result155[2]^and_result155[3]^and_result155[4]^and_result155[5]^and_result155[6]^and_result155[7]^and_result155[8]^and_result155[9]^and_result155[10]^and_result155[11]^and_result155[12]^and_result155[13]^and_result155[14]^and_result155[15]^and_result155[16]^and_result155[17]^and_result155[18]^and_result155[19]^and_result155[20]^and_result155[21]^and_result155[22]^and_result155[23]^and_result155[24]^and_result155[25]^and_result155[26]^and_result155[27]^and_result155[28]^and_result155[29]^and_result155[30]^and_result155[31]^and_result155[32]^and_result155[33]^and_result155[34]^and_result155[35]^and_result155[36]^and_result155[37]^and_result155[38]^and_result155[39]^and_result155[40]^and_result155[41]^and_result155[42]^and_result155[43]^and_result155[44]^and_result155[45]^and_result155[46]^and_result155[47]^and_result155[48]^and_result155[49]^and_result155[50]^and_result155[51]^and_result155[52]^and_result155[53]^and_result155[54]^and_result155[55]^and_result155[56]^and_result155[57]^and_result155[58]^and_result155[59]^and_result155[60]^and_result155[61]^and_result155[62]^and_result155[63]^and_result155[64]^and_result155[65]^and_result155[66]^and_result155[67]^and_result155[68]^and_result155[69]^and_result155[70]^and_result155[71]^and_result155[72]^and_result155[73]^and_result155[74]^and_result155[75]^and_result155[76]^and_result155[77]^and_result155[78]^and_result155[79]^and_result155[80]^and_result155[81]^and_result155[82]^and_result155[83]^and_result155[84]^and_result155[85]^and_result155[86]^and_result155[87]^and_result155[88]^and_result155[89]^and_result155[90]^and_result155[91]^and_result155[92]^and_result155[93]^and_result155[94]^and_result155[95]^and_result155[96]^and_result155[97]^and_result155[98]^and_result155[99]^and_result155[100]^and_result155[101]^and_result155[102]^and_result155[103]^and_result155[104]^and_result155[105]^and_result155[106]^and_result155[107]^and_result155[108]^and_result155[109]^and_result155[110]^and_result155[111]^and_result155[112]^and_result155[113]^and_result155[114]^and_result155[115]^and_result155[116]^and_result155[117]^and_result155[118]^and_result155[119]^and_result155[120]^and_result155[121]^and_result155[122]^and_result155[123]^and_result155[124]^and_result155[125]^and_result155[126]^and_result155[127]^and_result155[128]^and_result155[129]^and_result155[130]^and_result155[131]^and_result155[132]^and_result155[133]^and_result155[134]^and_result155[135]^and_result155[136]^and_result155[137]^and_result155[138]^and_result155[139]^and_result155[140]^and_result155[141]^and_result155[142]^and_result155[143]^and_result155[144]^and_result155[145]^and_result155[146]^and_result155[147]^and_result155[148]^and_result155[149]^and_result155[150]^and_result155[151]^and_result155[152]^and_result155[153]^and_result155[154]^and_result155[155]^and_result155[156]^and_result155[157]^and_result155[158]^and_result155[159]^and_result155[160]^and_result155[161]^and_result155[162]^and_result155[163]^and_result155[164]^and_result155[165]^and_result155[166]^and_result155[167]^and_result155[168]^and_result155[169]^and_result155[170]^and_result155[171]^and_result155[172]^and_result155[173]^and_result155[174]^and_result155[175]^and_result155[176]^and_result155[177]^and_result155[178]^and_result155[179]^and_result155[180]^and_result155[181]^and_result155[182]^and_result155[183]^and_result155[184]^and_result155[185]^and_result155[186]^and_result155[187]^and_result155[188]^and_result155[189]^and_result155[190]^and_result155[191]^and_result155[192]^and_result155[193]^and_result155[194]^and_result155[195]^and_result155[196]^and_result155[197]^and_result155[198]^and_result155[199]^and_result155[200]^and_result155[201]^and_result155[202]^and_result155[203]^and_result155[204]^and_result155[205]^and_result155[206]^and_result155[207]^and_result155[208]^and_result155[209]^and_result155[210]^and_result155[211]^and_result155[212]^and_result155[213]^and_result155[214]^and_result155[215]^and_result155[216]^and_result155[217]^and_result155[218]^and_result155[219]^and_result155[220]^and_result155[221]^and_result155[222]^and_result155[223]^and_result155[224]^and_result155[225]^and_result155[226]^and_result155[227]^and_result155[228]^and_result155[229]^and_result155[230]^and_result155[231]^and_result155[232]^and_result155[233]^and_result155[234]^and_result155[235]^and_result155[236]^and_result155[237]^and_result155[238]^and_result155[239]^and_result155[240]^and_result155[241]^and_result155[242]^and_result155[243]^and_result155[244]^and_result155[245]^and_result155[246]^and_result155[247]^and_result155[248]^and_result155[249]^and_result155[250]^and_result155[251]^and_result155[252]^and_result155[253]^and_result155[254];
assign key[156]=and_result156[0]^and_result156[1]^and_result156[2]^and_result156[3]^and_result156[4]^and_result156[5]^and_result156[6]^and_result156[7]^and_result156[8]^and_result156[9]^and_result156[10]^and_result156[11]^and_result156[12]^and_result156[13]^and_result156[14]^and_result156[15]^and_result156[16]^and_result156[17]^and_result156[18]^and_result156[19]^and_result156[20]^and_result156[21]^and_result156[22]^and_result156[23]^and_result156[24]^and_result156[25]^and_result156[26]^and_result156[27]^and_result156[28]^and_result156[29]^and_result156[30]^and_result156[31]^and_result156[32]^and_result156[33]^and_result156[34]^and_result156[35]^and_result156[36]^and_result156[37]^and_result156[38]^and_result156[39]^and_result156[40]^and_result156[41]^and_result156[42]^and_result156[43]^and_result156[44]^and_result156[45]^and_result156[46]^and_result156[47]^and_result156[48]^and_result156[49]^and_result156[50]^and_result156[51]^and_result156[52]^and_result156[53]^and_result156[54]^and_result156[55]^and_result156[56]^and_result156[57]^and_result156[58]^and_result156[59]^and_result156[60]^and_result156[61]^and_result156[62]^and_result156[63]^and_result156[64]^and_result156[65]^and_result156[66]^and_result156[67]^and_result156[68]^and_result156[69]^and_result156[70]^and_result156[71]^and_result156[72]^and_result156[73]^and_result156[74]^and_result156[75]^and_result156[76]^and_result156[77]^and_result156[78]^and_result156[79]^and_result156[80]^and_result156[81]^and_result156[82]^and_result156[83]^and_result156[84]^and_result156[85]^and_result156[86]^and_result156[87]^and_result156[88]^and_result156[89]^and_result156[90]^and_result156[91]^and_result156[92]^and_result156[93]^and_result156[94]^and_result156[95]^and_result156[96]^and_result156[97]^and_result156[98]^and_result156[99]^and_result156[100]^and_result156[101]^and_result156[102]^and_result156[103]^and_result156[104]^and_result156[105]^and_result156[106]^and_result156[107]^and_result156[108]^and_result156[109]^and_result156[110]^and_result156[111]^and_result156[112]^and_result156[113]^and_result156[114]^and_result156[115]^and_result156[116]^and_result156[117]^and_result156[118]^and_result156[119]^and_result156[120]^and_result156[121]^and_result156[122]^and_result156[123]^and_result156[124]^and_result156[125]^and_result156[126]^and_result156[127]^and_result156[128]^and_result156[129]^and_result156[130]^and_result156[131]^and_result156[132]^and_result156[133]^and_result156[134]^and_result156[135]^and_result156[136]^and_result156[137]^and_result156[138]^and_result156[139]^and_result156[140]^and_result156[141]^and_result156[142]^and_result156[143]^and_result156[144]^and_result156[145]^and_result156[146]^and_result156[147]^and_result156[148]^and_result156[149]^and_result156[150]^and_result156[151]^and_result156[152]^and_result156[153]^and_result156[154]^and_result156[155]^and_result156[156]^and_result156[157]^and_result156[158]^and_result156[159]^and_result156[160]^and_result156[161]^and_result156[162]^and_result156[163]^and_result156[164]^and_result156[165]^and_result156[166]^and_result156[167]^and_result156[168]^and_result156[169]^and_result156[170]^and_result156[171]^and_result156[172]^and_result156[173]^and_result156[174]^and_result156[175]^and_result156[176]^and_result156[177]^and_result156[178]^and_result156[179]^and_result156[180]^and_result156[181]^and_result156[182]^and_result156[183]^and_result156[184]^and_result156[185]^and_result156[186]^and_result156[187]^and_result156[188]^and_result156[189]^and_result156[190]^and_result156[191]^and_result156[192]^and_result156[193]^and_result156[194]^and_result156[195]^and_result156[196]^and_result156[197]^and_result156[198]^and_result156[199]^and_result156[200]^and_result156[201]^and_result156[202]^and_result156[203]^and_result156[204]^and_result156[205]^and_result156[206]^and_result156[207]^and_result156[208]^and_result156[209]^and_result156[210]^and_result156[211]^and_result156[212]^and_result156[213]^and_result156[214]^and_result156[215]^and_result156[216]^and_result156[217]^and_result156[218]^and_result156[219]^and_result156[220]^and_result156[221]^and_result156[222]^and_result156[223]^and_result156[224]^and_result156[225]^and_result156[226]^and_result156[227]^and_result156[228]^and_result156[229]^and_result156[230]^and_result156[231]^and_result156[232]^and_result156[233]^and_result156[234]^and_result156[235]^and_result156[236]^and_result156[237]^and_result156[238]^and_result156[239]^and_result156[240]^and_result156[241]^and_result156[242]^and_result156[243]^and_result156[244]^and_result156[245]^and_result156[246]^and_result156[247]^and_result156[248]^and_result156[249]^and_result156[250]^and_result156[251]^and_result156[252]^and_result156[253]^and_result156[254];
assign key[157]=and_result157[0]^and_result157[1]^and_result157[2]^and_result157[3]^and_result157[4]^and_result157[5]^and_result157[6]^and_result157[7]^and_result157[8]^and_result157[9]^and_result157[10]^and_result157[11]^and_result157[12]^and_result157[13]^and_result157[14]^and_result157[15]^and_result157[16]^and_result157[17]^and_result157[18]^and_result157[19]^and_result157[20]^and_result157[21]^and_result157[22]^and_result157[23]^and_result157[24]^and_result157[25]^and_result157[26]^and_result157[27]^and_result157[28]^and_result157[29]^and_result157[30]^and_result157[31]^and_result157[32]^and_result157[33]^and_result157[34]^and_result157[35]^and_result157[36]^and_result157[37]^and_result157[38]^and_result157[39]^and_result157[40]^and_result157[41]^and_result157[42]^and_result157[43]^and_result157[44]^and_result157[45]^and_result157[46]^and_result157[47]^and_result157[48]^and_result157[49]^and_result157[50]^and_result157[51]^and_result157[52]^and_result157[53]^and_result157[54]^and_result157[55]^and_result157[56]^and_result157[57]^and_result157[58]^and_result157[59]^and_result157[60]^and_result157[61]^and_result157[62]^and_result157[63]^and_result157[64]^and_result157[65]^and_result157[66]^and_result157[67]^and_result157[68]^and_result157[69]^and_result157[70]^and_result157[71]^and_result157[72]^and_result157[73]^and_result157[74]^and_result157[75]^and_result157[76]^and_result157[77]^and_result157[78]^and_result157[79]^and_result157[80]^and_result157[81]^and_result157[82]^and_result157[83]^and_result157[84]^and_result157[85]^and_result157[86]^and_result157[87]^and_result157[88]^and_result157[89]^and_result157[90]^and_result157[91]^and_result157[92]^and_result157[93]^and_result157[94]^and_result157[95]^and_result157[96]^and_result157[97]^and_result157[98]^and_result157[99]^and_result157[100]^and_result157[101]^and_result157[102]^and_result157[103]^and_result157[104]^and_result157[105]^and_result157[106]^and_result157[107]^and_result157[108]^and_result157[109]^and_result157[110]^and_result157[111]^and_result157[112]^and_result157[113]^and_result157[114]^and_result157[115]^and_result157[116]^and_result157[117]^and_result157[118]^and_result157[119]^and_result157[120]^and_result157[121]^and_result157[122]^and_result157[123]^and_result157[124]^and_result157[125]^and_result157[126]^and_result157[127]^and_result157[128]^and_result157[129]^and_result157[130]^and_result157[131]^and_result157[132]^and_result157[133]^and_result157[134]^and_result157[135]^and_result157[136]^and_result157[137]^and_result157[138]^and_result157[139]^and_result157[140]^and_result157[141]^and_result157[142]^and_result157[143]^and_result157[144]^and_result157[145]^and_result157[146]^and_result157[147]^and_result157[148]^and_result157[149]^and_result157[150]^and_result157[151]^and_result157[152]^and_result157[153]^and_result157[154]^and_result157[155]^and_result157[156]^and_result157[157]^and_result157[158]^and_result157[159]^and_result157[160]^and_result157[161]^and_result157[162]^and_result157[163]^and_result157[164]^and_result157[165]^and_result157[166]^and_result157[167]^and_result157[168]^and_result157[169]^and_result157[170]^and_result157[171]^and_result157[172]^and_result157[173]^and_result157[174]^and_result157[175]^and_result157[176]^and_result157[177]^and_result157[178]^and_result157[179]^and_result157[180]^and_result157[181]^and_result157[182]^and_result157[183]^and_result157[184]^and_result157[185]^and_result157[186]^and_result157[187]^and_result157[188]^and_result157[189]^and_result157[190]^and_result157[191]^and_result157[192]^and_result157[193]^and_result157[194]^and_result157[195]^and_result157[196]^and_result157[197]^and_result157[198]^and_result157[199]^and_result157[200]^and_result157[201]^and_result157[202]^and_result157[203]^and_result157[204]^and_result157[205]^and_result157[206]^and_result157[207]^and_result157[208]^and_result157[209]^and_result157[210]^and_result157[211]^and_result157[212]^and_result157[213]^and_result157[214]^and_result157[215]^and_result157[216]^and_result157[217]^and_result157[218]^and_result157[219]^and_result157[220]^and_result157[221]^and_result157[222]^and_result157[223]^and_result157[224]^and_result157[225]^and_result157[226]^and_result157[227]^and_result157[228]^and_result157[229]^and_result157[230]^and_result157[231]^and_result157[232]^and_result157[233]^and_result157[234]^and_result157[235]^and_result157[236]^and_result157[237]^and_result157[238]^and_result157[239]^and_result157[240]^and_result157[241]^and_result157[242]^and_result157[243]^and_result157[244]^and_result157[245]^and_result157[246]^and_result157[247]^and_result157[248]^and_result157[249]^and_result157[250]^and_result157[251]^and_result157[252]^and_result157[253]^and_result157[254];
assign key[158]=and_result158[0]^and_result158[1]^and_result158[2]^and_result158[3]^and_result158[4]^and_result158[5]^and_result158[6]^and_result158[7]^and_result158[8]^and_result158[9]^and_result158[10]^and_result158[11]^and_result158[12]^and_result158[13]^and_result158[14]^and_result158[15]^and_result158[16]^and_result158[17]^and_result158[18]^and_result158[19]^and_result158[20]^and_result158[21]^and_result158[22]^and_result158[23]^and_result158[24]^and_result158[25]^and_result158[26]^and_result158[27]^and_result158[28]^and_result158[29]^and_result158[30]^and_result158[31]^and_result158[32]^and_result158[33]^and_result158[34]^and_result158[35]^and_result158[36]^and_result158[37]^and_result158[38]^and_result158[39]^and_result158[40]^and_result158[41]^and_result158[42]^and_result158[43]^and_result158[44]^and_result158[45]^and_result158[46]^and_result158[47]^and_result158[48]^and_result158[49]^and_result158[50]^and_result158[51]^and_result158[52]^and_result158[53]^and_result158[54]^and_result158[55]^and_result158[56]^and_result158[57]^and_result158[58]^and_result158[59]^and_result158[60]^and_result158[61]^and_result158[62]^and_result158[63]^and_result158[64]^and_result158[65]^and_result158[66]^and_result158[67]^and_result158[68]^and_result158[69]^and_result158[70]^and_result158[71]^and_result158[72]^and_result158[73]^and_result158[74]^and_result158[75]^and_result158[76]^and_result158[77]^and_result158[78]^and_result158[79]^and_result158[80]^and_result158[81]^and_result158[82]^and_result158[83]^and_result158[84]^and_result158[85]^and_result158[86]^and_result158[87]^and_result158[88]^and_result158[89]^and_result158[90]^and_result158[91]^and_result158[92]^and_result158[93]^and_result158[94]^and_result158[95]^and_result158[96]^and_result158[97]^and_result158[98]^and_result158[99]^and_result158[100]^and_result158[101]^and_result158[102]^and_result158[103]^and_result158[104]^and_result158[105]^and_result158[106]^and_result158[107]^and_result158[108]^and_result158[109]^and_result158[110]^and_result158[111]^and_result158[112]^and_result158[113]^and_result158[114]^and_result158[115]^and_result158[116]^and_result158[117]^and_result158[118]^and_result158[119]^and_result158[120]^and_result158[121]^and_result158[122]^and_result158[123]^and_result158[124]^and_result158[125]^and_result158[126]^and_result158[127]^and_result158[128]^and_result158[129]^and_result158[130]^and_result158[131]^and_result158[132]^and_result158[133]^and_result158[134]^and_result158[135]^and_result158[136]^and_result158[137]^and_result158[138]^and_result158[139]^and_result158[140]^and_result158[141]^and_result158[142]^and_result158[143]^and_result158[144]^and_result158[145]^and_result158[146]^and_result158[147]^and_result158[148]^and_result158[149]^and_result158[150]^and_result158[151]^and_result158[152]^and_result158[153]^and_result158[154]^and_result158[155]^and_result158[156]^and_result158[157]^and_result158[158]^and_result158[159]^and_result158[160]^and_result158[161]^and_result158[162]^and_result158[163]^and_result158[164]^and_result158[165]^and_result158[166]^and_result158[167]^and_result158[168]^and_result158[169]^and_result158[170]^and_result158[171]^and_result158[172]^and_result158[173]^and_result158[174]^and_result158[175]^and_result158[176]^and_result158[177]^and_result158[178]^and_result158[179]^and_result158[180]^and_result158[181]^and_result158[182]^and_result158[183]^and_result158[184]^and_result158[185]^and_result158[186]^and_result158[187]^and_result158[188]^and_result158[189]^and_result158[190]^and_result158[191]^and_result158[192]^and_result158[193]^and_result158[194]^and_result158[195]^and_result158[196]^and_result158[197]^and_result158[198]^and_result158[199]^and_result158[200]^and_result158[201]^and_result158[202]^and_result158[203]^and_result158[204]^and_result158[205]^and_result158[206]^and_result158[207]^and_result158[208]^and_result158[209]^and_result158[210]^and_result158[211]^and_result158[212]^and_result158[213]^and_result158[214]^and_result158[215]^and_result158[216]^and_result158[217]^and_result158[218]^and_result158[219]^and_result158[220]^and_result158[221]^and_result158[222]^and_result158[223]^and_result158[224]^and_result158[225]^and_result158[226]^and_result158[227]^and_result158[228]^and_result158[229]^and_result158[230]^and_result158[231]^and_result158[232]^and_result158[233]^and_result158[234]^and_result158[235]^and_result158[236]^and_result158[237]^and_result158[238]^and_result158[239]^and_result158[240]^and_result158[241]^and_result158[242]^and_result158[243]^and_result158[244]^and_result158[245]^and_result158[246]^and_result158[247]^and_result158[248]^and_result158[249]^and_result158[250]^and_result158[251]^and_result158[252]^and_result158[253]^and_result158[254];
assign key[159]=and_result159[0]^and_result159[1]^and_result159[2]^and_result159[3]^and_result159[4]^and_result159[5]^and_result159[6]^and_result159[7]^and_result159[8]^and_result159[9]^and_result159[10]^and_result159[11]^and_result159[12]^and_result159[13]^and_result159[14]^and_result159[15]^and_result159[16]^and_result159[17]^and_result159[18]^and_result159[19]^and_result159[20]^and_result159[21]^and_result159[22]^and_result159[23]^and_result159[24]^and_result159[25]^and_result159[26]^and_result159[27]^and_result159[28]^and_result159[29]^and_result159[30]^and_result159[31]^and_result159[32]^and_result159[33]^and_result159[34]^and_result159[35]^and_result159[36]^and_result159[37]^and_result159[38]^and_result159[39]^and_result159[40]^and_result159[41]^and_result159[42]^and_result159[43]^and_result159[44]^and_result159[45]^and_result159[46]^and_result159[47]^and_result159[48]^and_result159[49]^and_result159[50]^and_result159[51]^and_result159[52]^and_result159[53]^and_result159[54]^and_result159[55]^and_result159[56]^and_result159[57]^and_result159[58]^and_result159[59]^and_result159[60]^and_result159[61]^and_result159[62]^and_result159[63]^and_result159[64]^and_result159[65]^and_result159[66]^and_result159[67]^and_result159[68]^and_result159[69]^and_result159[70]^and_result159[71]^and_result159[72]^and_result159[73]^and_result159[74]^and_result159[75]^and_result159[76]^and_result159[77]^and_result159[78]^and_result159[79]^and_result159[80]^and_result159[81]^and_result159[82]^and_result159[83]^and_result159[84]^and_result159[85]^and_result159[86]^and_result159[87]^and_result159[88]^and_result159[89]^and_result159[90]^and_result159[91]^and_result159[92]^and_result159[93]^and_result159[94]^and_result159[95]^and_result159[96]^and_result159[97]^and_result159[98]^and_result159[99]^and_result159[100]^and_result159[101]^and_result159[102]^and_result159[103]^and_result159[104]^and_result159[105]^and_result159[106]^and_result159[107]^and_result159[108]^and_result159[109]^and_result159[110]^and_result159[111]^and_result159[112]^and_result159[113]^and_result159[114]^and_result159[115]^and_result159[116]^and_result159[117]^and_result159[118]^and_result159[119]^and_result159[120]^and_result159[121]^and_result159[122]^and_result159[123]^and_result159[124]^and_result159[125]^and_result159[126]^and_result159[127]^and_result159[128]^and_result159[129]^and_result159[130]^and_result159[131]^and_result159[132]^and_result159[133]^and_result159[134]^and_result159[135]^and_result159[136]^and_result159[137]^and_result159[138]^and_result159[139]^and_result159[140]^and_result159[141]^and_result159[142]^and_result159[143]^and_result159[144]^and_result159[145]^and_result159[146]^and_result159[147]^and_result159[148]^and_result159[149]^and_result159[150]^and_result159[151]^and_result159[152]^and_result159[153]^and_result159[154]^and_result159[155]^and_result159[156]^and_result159[157]^and_result159[158]^and_result159[159]^and_result159[160]^and_result159[161]^and_result159[162]^and_result159[163]^and_result159[164]^and_result159[165]^and_result159[166]^and_result159[167]^and_result159[168]^and_result159[169]^and_result159[170]^and_result159[171]^and_result159[172]^and_result159[173]^and_result159[174]^and_result159[175]^and_result159[176]^and_result159[177]^and_result159[178]^and_result159[179]^and_result159[180]^and_result159[181]^and_result159[182]^and_result159[183]^and_result159[184]^and_result159[185]^and_result159[186]^and_result159[187]^and_result159[188]^and_result159[189]^and_result159[190]^and_result159[191]^and_result159[192]^and_result159[193]^and_result159[194]^and_result159[195]^and_result159[196]^and_result159[197]^and_result159[198]^and_result159[199]^and_result159[200]^and_result159[201]^and_result159[202]^and_result159[203]^and_result159[204]^and_result159[205]^and_result159[206]^and_result159[207]^and_result159[208]^and_result159[209]^and_result159[210]^and_result159[211]^and_result159[212]^and_result159[213]^and_result159[214]^and_result159[215]^and_result159[216]^and_result159[217]^and_result159[218]^and_result159[219]^and_result159[220]^and_result159[221]^and_result159[222]^and_result159[223]^and_result159[224]^and_result159[225]^and_result159[226]^and_result159[227]^and_result159[228]^and_result159[229]^and_result159[230]^and_result159[231]^and_result159[232]^and_result159[233]^and_result159[234]^and_result159[235]^and_result159[236]^and_result159[237]^and_result159[238]^and_result159[239]^and_result159[240]^and_result159[241]^and_result159[242]^and_result159[243]^and_result159[244]^and_result159[245]^and_result159[246]^and_result159[247]^and_result159[248]^and_result159[249]^and_result159[250]^and_result159[251]^and_result159[252]^and_result159[253]^and_result159[254];
assign key[160]=and_result160[0]^and_result160[1]^and_result160[2]^and_result160[3]^and_result160[4]^and_result160[5]^and_result160[6]^and_result160[7]^and_result160[8]^and_result160[9]^and_result160[10]^and_result160[11]^and_result160[12]^and_result160[13]^and_result160[14]^and_result160[15]^and_result160[16]^and_result160[17]^and_result160[18]^and_result160[19]^and_result160[20]^and_result160[21]^and_result160[22]^and_result160[23]^and_result160[24]^and_result160[25]^and_result160[26]^and_result160[27]^and_result160[28]^and_result160[29]^and_result160[30]^and_result160[31]^and_result160[32]^and_result160[33]^and_result160[34]^and_result160[35]^and_result160[36]^and_result160[37]^and_result160[38]^and_result160[39]^and_result160[40]^and_result160[41]^and_result160[42]^and_result160[43]^and_result160[44]^and_result160[45]^and_result160[46]^and_result160[47]^and_result160[48]^and_result160[49]^and_result160[50]^and_result160[51]^and_result160[52]^and_result160[53]^and_result160[54]^and_result160[55]^and_result160[56]^and_result160[57]^and_result160[58]^and_result160[59]^and_result160[60]^and_result160[61]^and_result160[62]^and_result160[63]^and_result160[64]^and_result160[65]^and_result160[66]^and_result160[67]^and_result160[68]^and_result160[69]^and_result160[70]^and_result160[71]^and_result160[72]^and_result160[73]^and_result160[74]^and_result160[75]^and_result160[76]^and_result160[77]^and_result160[78]^and_result160[79]^and_result160[80]^and_result160[81]^and_result160[82]^and_result160[83]^and_result160[84]^and_result160[85]^and_result160[86]^and_result160[87]^and_result160[88]^and_result160[89]^and_result160[90]^and_result160[91]^and_result160[92]^and_result160[93]^and_result160[94]^and_result160[95]^and_result160[96]^and_result160[97]^and_result160[98]^and_result160[99]^and_result160[100]^and_result160[101]^and_result160[102]^and_result160[103]^and_result160[104]^and_result160[105]^and_result160[106]^and_result160[107]^and_result160[108]^and_result160[109]^and_result160[110]^and_result160[111]^and_result160[112]^and_result160[113]^and_result160[114]^and_result160[115]^and_result160[116]^and_result160[117]^and_result160[118]^and_result160[119]^and_result160[120]^and_result160[121]^and_result160[122]^and_result160[123]^and_result160[124]^and_result160[125]^and_result160[126]^and_result160[127]^and_result160[128]^and_result160[129]^and_result160[130]^and_result160[131]^and_result160[132]^and_result160[133]^and_result160[134]^and_result160[135]^and_result160[136]^and_result160[137]^and_result160[138]^and_result160[139]^and_result160[140]^and_result160[141]^and_result160[142]^and_result160[143]^and_result160[144]^and_result160[145]^and_result160[146]^and_result160[147]^and_result160[148]^and_result160[149]^and_result160[150]^and_result160[151]^and_result160[152]^and_result160[153]^and_result160[154]^and_result160[155]^and_result160[156]^and_result160[157]^and_result160[158]^and_result160[159]^and_result160[160]^and_result160[161]^and_result160[162]^and_result160[163]^and_result160[164]^and_result160[165]^and_result160[166]^and_result160[167]^and_result160[168]^and_result160[169]^and_result160[170]^and_result160[171]^and_result160[172]^and_result160[173]^and_result160[174]^and_result160[175]^and_result160[176]^and_result160[177]^and_result160[178]^and_result160[179]^and_result160[180]^and_result160[181]^and_result160[182]^and_result160[183]^and_result160[184]^and_result160[185]^and_result160[186]^and_result160[187]^and_result160[188]^and_result160[189]^and_result160[190]^and_result160[191]^and_result160[192]^and_result160[193]^and_result160[194]^and_result160[195]^and_result160[196]^and_result160[197]^and_result160[198]^and_result160[199]^and_result160[200]^and_result160[201]^and_result160[202]^and_result160[203]^and_result160[204]^and_result160[205]^and_result160[206]^and_result160[207]^and_result160[208]^and_result160[209]^and_result160[210]^and_result160[211]^and_result160[212]^and_result160[213]^and_result160[214]^and_result160[215]^and_result160[216]^and_result160[217]^and_result160[218]^and_result160[219]^and_result160[220]^and_result160[221]^and_result160[222]^and_result160[223]^and_result160[224]^and_result160[225]^and_result160[226]^and_result160[227]^and_result160[228]^and_result160[229]^and_result160[230]^and_result160[231]^and_result160[232]^and_result160[233]^and_result160[234]^and_result160[235]^and_result160[236]^and_result160[237]^and_result160[238]^and_result160[239]^and_result160[240]^and_result160[241]^and_result160[242]^and_result160[243]^and_result160[244]^and_result160[245]^and_result160[246]^and_result160[247]^and_result160[248]^and_result160[249]^and_result160[250]^and_result160[251]^and_result160[252]^and_result160[253]^and_result160[254];
assign key[161]=and_result161[0]^and_result161[1]^and_result161[2]^and_result161[3]^and_result161[4]^and_result161[5]^and_result161[6]^and_result161[7]^and_result161[8]^and_result161[9]^and_result161[10]^and_result161[11]^and_result161[12]^and_result161[13]^and_result161[14]^and_result161[15]^and_result161[16]^and_result161[17]^and_result161[18]^and_result161[19]^and_result161[20]^and_result161[21]^and_result161[22]^and_result161[23]^and_result161[24]^and_result161[25]^and_result161[26]^and_result161[27]^and_result161[28]^and_result161[29]^and_result161[30]^and_result161[31]^and_result161[32]^and_result161[33]^and_result161[34]^and_result161[35]^and_result161[36]^and_result161[37]^and_result161[38]^and_result161[39]^and_result161[40]^and_result161[41]^and_result161[42]^and_result161[43]^and_result161[44]^and_result161[45]^and_result161[46]^and_result161[47]^and_result161[48]^and_result161[49]^and_result161[50]^and_result161[51]^and_result161[52]^and_result161[53]^and_result161[54]^and_result161[55]^and_result161[56]^and_result161[57]^and_result161[58]^and_result161[59]^and_result161[60]^and_result161[61]^and_result161[62]^and_result161[63]^and_result161[64]^and_result161[65]^and_result161[66]^and_result161[67]^and_result161[68]^and_result161[69]^and_result161[70]^and_result161[71]^and_result161[72]^and_result161[73]^and_result161[74]^and_result161[75]^and_result161[76]^and_result161[77]^and_result161[78]^and_result161[79]^and_result161[80]^and_result161[81]^and_result161[82]^and_result161[83]^and_result161[84]^and_result161[85]^and_result161[86]^and_result161[87]^and_result161[88]^and_result161[89]^and_result161[90]^and_result161[91]^and_result161[92]^and_result161[93]^and_result161[94]^and_result161[95]^and_result161[96]^and_result161[97]^and_result161[98]^and_result161[99]^and_result161[100]^and_result161[101]^and_result161[102]^and_result161[103]^and_result161[104]^and_result161[105]^and_result161[106]^and_result161[107]^and_result161[108]^and_result161[109]^and_result161[110]^and_result161[111]^and_result161[112]^and_result161[113]^and_result161[114]^and_result161[115]^and_result161[116]^and_result161[117]^and_result161[118]^and_result161[119]^and_result161[120]^and_result161[121]^and_result161[122]^and_result161[123]^and_result161[124]^and_result161[125]^and_result161[126]^and_result161[127]^and_result161[128]^and_result161[129]^and_result161[130]^and_result161[131]^and_result161[132]^and_result161[133]^and_result161[134]^and_result161[135]^and_result161[136]^and_result161[137]^and_result161[138]^and_result161[139]^and_result161[140]^and_result161[141]^and_result161[142]^and_result161[143]^and_result161[144]^and_result161[145]^and_result161[146]^and_result161[147]^and_result161[148]^and_result161[149]^and_result161[150]^and_result161[151]^and_result161[152]^and_result161[153]^and_result161[154]^and_result161[155]^and_result161[156]^and_result161[157]^and_result161[158]^and_result161[159]^and_result161[160]^and_result161[161]^and_result161[162]^and_result161[163]^and_result161[164]^and_result161[165]^and_result161[166]^and_result161[167]^and_result161[168]^and_result161[169]^and_result161[170]^and_result161[171]^and_result161[172]^and_result161[173]^and_result161[174]^and_result161[175]^and_result161[176]^and_result161[177]^and_result161[178]^and_result161[179]^and_result161[180]^and_result161[181]^and_result161[182]^and_result161[183]^and_result161[184]^and_result161[185]^and_result161[186]^and_result161[187]^and_result161[188]^and_result161[189]^and_result161[190]^and_result161[191]^and_result161[192]^and_result161[193]^and_result161[194]^and_result161[195]^and_result161[196]^and_result161[197]^and_result161[198]^and_result161[199]^and_result161[200]^and_result161[201]^and_result161[202]^and_result161[203]^and_result161[204]^and_result161[205]^and_result161[206]^and_result161[207]^and_result161[208]^and_result161[209]^and_result161[210]^and_result161[211]^and_result161[212]^and_result161[213]^and_result161[214]^and_result161[215]^and_result161[216]^and_result161[217]^and_result161[218]^and_result161[219]^and_result161[220]^and_result161[221]^and_result161[222]^and_result161[223]^and_result161[224]^and_result161[225]^and_result161[226]^and_result161[227]^and_result161[228]^and_result161[229]^and_result161[230]^and_result161[231]^and_result161[232]^and_result161[233]^and_result161[234]^and_result161[235]^and_result161[236]^and_result161[237]^and_result161[238]^and_result161[239]^and_result161[240]^and_result161[241]^and_result161[242]^and_result161[243]^and_result161[244]^and_result161[245]^and_result161[246]^and_result161[247]^and_result161[248]^and_result161[249]^and_result161[250]^and_result161[251]^and_result161[252]^and_result161[253]^and_result161[254];
assign key[162]=and_result162[0]^and_result162[1]^and_result162[2]^and_result162[3]^and_result162[4]^and_result162[5]^and_result162[6]^and_result162[7]^and_result162[8]^and_result162[9]^and_result162[10]^and_result162[11]^and_result162[12]^and_result162[13]^and_result162[14]^and_result162[15]^and_result162[16]^and_result162[17]^and_result162[18]^and_result162[19]^and_result162[20]^and_result162[21]^and_result162[22]^and_result162[23]^and_result162[24]^and_result162[25]^and_result162[26]^and_result162[27]^and_result162[28]^and_result162[29]^and_result162[30]^and_result162[31]^and_result162[32]^and_result162[33]^and_result162[34]^and_result162[35]^and_result162[36]^and_result162[37]^and_result162[38]^and_result162[39]^and_result162[40]^and_result162[41]^and_result162[42]^and_result162[43]^and_result162[44]^and_result162[45]^and_result162[46]^and_result162[47]^and_result162[48]^and_result162[49]^and_result162[50]^and_result162[51]^and_result162[52]^and_result162[53]^and_result162[54]^and_result162[55]^and_result162[56]^and_result162[57]^and_result162[58]^and_result162[59]^and_result162[60]^and_result162[61]^and_result162[62]^and_result162[63]^and_result162[64]^and_result162[65]^and_result162[66]^and_result162[67]^and_result162[68]^and_result162[69]^and_result162[70]^and_result162[71]^and_result162[72]^and_result162[73]^and_result162[74]^and_result162[75]^and_result162[76]^and_result162[77]^and_result162[78]^and_result162[79]^and_result162[80]^and_result162[81]^and_result162[82]^and_result162[83]^and_result162[84]^and_result162[85]^and_result162[86]^and_result162[87]^and_result162[88]^and_result162[89]^and_result162[90]^and_result162[91]^and_result162[92]^and_result162[93]^and_result162[94]^and_result162[95]^and_result162[96]^and_result162[97]^and_result162[98]^and_result162[99]^and_result162[100]^and_result162[101]^and_result162[102]^and_result162[103]^and_result162[104]^and_result162[105]^and_result162[106]^and_result162[107]^and_result162[108]^and_result162[109]^and_result162[110]^and_result162[111]^and_result162[112]^and_result162[113]^and_result162[114]^and_result162[115]^and_result162[116]^and_result162[117]^and_result162[118]^and_result162[119]^and_result162[120]^and_result162[121]^and_result162[122]^and_result162[123]^and_result162[124]^and_result162[125]^and_result162[126]^and_result162[127]^and_result162[128]^and_result162[129]^and_result162[130]^and_result162[131]^and_result162[132]^and_result162[133]^and_result162[134]^and_result162[135]^and_result162[136]^and_result162[137]^and_result162[138]^and_result162[139]^and_result162[140]^and_result162[141]^and_result162[142]^and_result162[143]^and_result162[144]^and_result162[145]^and_result162[146]^and_result162[147]^and_result162[148]^and_result162[149]^and_result162[150]^and_result162[151]^and_result162[152]^and_result162[153]^and_result162[154]^and_result162[155]^and_result162[156]^and_result162[157]^and_result162[158]^and_result162[159]^and_result162[160]^and_result162[161]^and_result162[162]^and_result162[163]^and_result162[164]^and_result162[165]^and_result162[166]^and_result162[167]^and_result162[168]^and_result162[169]^and_result162[170]^and_result162[171]^and_result162[172]^and_result162[173]^and_result162[174]^and_result162[175]^and_result162[176]^and_result162[177]^and_result162[178]^and_result162[179]^and_result162[180]^and_result162[181]^and_result162[182]^and_result162[183]^and_result162[184]^and_result162[185]^and_result162[186]^and_result162[187]^and_result162[188]^and_result162[189]^and_result162[190]^and_result162[191]^and_result162[192]^and_result162[193]^and_result162[194]^and_result162[195]^and_result162[196]^and_result162[197]^and_result162[198]^and_result162[199]^and_result162[200]^and_result162[201]^and_result162[202]^and_result162[203]^and_result162[204]^and_result162[205]^and_result162[206]^and_result162[207]^and_result162[208]^and_result162[209]^and_result162[210]^and_result162[211]^and_result162[212]^and_result162[213]^and_result162[214]^and_result162[215]^and_result162[216]^and_result162[217]^and_result162[218]^and_result162[219]^and_result162[220]^and_result162[221]^and_result162[222]^and_result162[223]^and_result162[224]^and_result162[225]^and_result162[226]^and_result162[227]^and_result162[228]^and_result162[229]^and_result162[230]^and_result162[231]^and_result162[232]^and_result162[233]^and_result162[234]^and_result162[235]^and_result162[236]^and_result162[237]^and_result162[238]^and_result162[239]^and_result162[240]^and_result162[241]^and_result162[242]^and_result162[243]^and_result162[244]^and_result162[245]^and_result162[246]^and_result162[247]^and_result162[248]^and_result162[249]^and_result162[250]^and_result162[251]^and_result162[252]^and_result162[253]^and_result162[254];
assign key[163]=and_result163[0]^and_result163[1]^and_result163[2]^and_result163[3]^and_result163[4]^and_result163[5]^and_result163[6]^and_result163[7]^and_result163[8]^and_result163[9]^and_result163[10]^and_result163[11]^and_result163[12]^and_result163[13]^and_result163[14]^and_result163[15]^and_result163[16]^and_result163[17]^and_result163[18]^and_result163[19]^and_result163[20]^and_result163[21]^and_result163[22]^and_result163[23]^and_result163[24]^and_result163[25]^and_result163[26]^and_result163[27]^and_result163[28]^and_result163[29]^and_result163[30]^and_result163[31]^and_result163[32]^and_result163[33]^and_result163[34]^and_result163[35]^and_result163[36]^and_result163[37]^and_result163[38]^and_result163[39]^and_result163[40]^and_result163[41]^and_result163[42]^and_result163[43]^and_result163[44]^and_result163[45]^and_result163[46]^and_result163[47]^and_result163[48]^and_result163[49]^and_result163[50]^and_result163[51]^and_result163[52]^and_result163[53]^and_result163[54]^and_result163[55]^and_result163[56]^and_result163[57]^and_result163[58]^and_result163[59]^and_result163[60]^and_result163[61]^and_result163[62]^and_result163[63]^and_result163[64]^and_result163[65]^and_result163[66]^and_result163[67]^and_result163[68]^and_result163[69]^and_result163[70]^and_result163[71]^and_result163[72]^and_result163[73]^and_result163[74]^and_result163[75]^and_result163[76]^and_result163[77]^and_result163[78]^and_result163[79]^and_result163[80]^and_result163[81]^and_result163[82]^and_result163[83]^and_result163[84]^and_result163[85]^and_result163[86]^and_result163[87]^and_result163[88]^and_result163[89]^and_result163[90]^and_result163[91]^and_result163[92]^and_result163[93]^and_result163[94]^and_result163[95]^and_result163[96]^and_result163[97]^and_result163[98]^and_result163[99]^and_result163[100]^and_result163[101]^and_result163[102]^and_result163[103]^and_result163[104]^and_result163[105]^and_result163[106]^and_result163[107]^and_result163[108]^and_result163[109]^and_result163[110]^and_result163[111]^and_result163[112]^and_result163[113]^and_result163[114]^and_result163[115]^and_result163[116]^and_result163[117]^and_result163[118]^and_result163[119]^and_result163[120]^and_result163[121]^and_result163[122]^and_result163[123]^and_result163[124]^and_result163[125]^and_result163[126]^and_result163[127]^and_result163[128]^and_result163[129]^and_result163[130]^and_result163[131]^and_result163[132]^and_result163[133]^and_result163[134]^and_result163[135]^and_result163[136]^and_result163[137]^and_result163[138]^and_result163[139]^and_result163[140]^and_result163[141]^and_result163[142]^and_result163[143]^and_result163[144]^and_result163[145]^and_result163[146]^and_result163[147]^and_result163[148]^and_result163[149]^and_result163[150]^and_result163[151]^and_result163[152]^and_result163[153]^and_result163[154]^and_result163[155]^and_result163[156]^and_result163[157]^and_result163[158]^and_result163[159]^and_result163[160]^and_result163[161]^and_result163[162]^and_result163[163]^and_result163[164]^and_result163[165]^and_result163[166]^and_result163[167]^and_result163[168]^and_result163[169]^and_result163[170]^and_result163[171]^and_result163[172]^and_result163[173]^and_result163[174]^and_result163[175]^and_result163[176]^and_result163[177]^and_result163[178]^and_result163[179]^and_result163[180]^and_result163[181]^and_result163[182]^and_result163[183]^and_result163[184]^and_result163[185]^and_result163[186]^and_result163[187]^and_result163[188]^and_result163[189]^and_result163[190]^and_result163[191]^and_result163[192]^and_result163[193]^and_result163[194]^and_result163[195]^and_result163[196]^and_result163[197]^and_result163[198]^and_result163[199]^and_result163[200]^and_result163[201]^and_result163[202]^and_result163[203]^and_result163[204]^and_result163[205]^and_result163[206]^and_result163[207]^and_result163[208]^and_result163[209]^and_result163[210]^and_result163[211]^and_result163[212]^and_result163[213]^and_result163[214]^and_result163[215]^and_result163[216]^and_result163[217]^and_result163[218]^and_result163[219]^and_result163[220]^and_result163[221]^and_result163[222]^and_result163[223]^and_result163[224]^and_result163[225]^and_result163[226]^and_result163[227]^and_result163[228]^and_result163[229]^and_result163[230]^and_result163[231]^and_result163[232]^and_result163[233]^and_result163[234]^and_result163[235]^and_result163[236]^and_result163[237]^and_result163[238]^and_result163[239]^and_result163[240]^and_result163[241]^and_result163[242]^and_result163[243]^and_result163[244]^and_result163[245]^and_result163[246]^and_result163[247]^and_result163[248]^and_result163[249]^and_result163[250]^and_result163[251]^and_result163[252]^and_result163[253]^and_result163[254];
assign key[164]=and_result164[0]^and_result164[1]^and_result164[2]^and_result164[3]^and_result164[4]^and_result164[5]^and_result164[6]^and_result164[7]^and_result164[8]^and_result164[9]^and_result164[10]^and_result164[11]^and_result164[12]^and_result164[13]^and_result164[14]^and_result164[15]^and_result164[16]^and_result164[17]^and_result164[18]^and_result164[19]^and_result164[20]^and_result164[21]^and_result164[22]^and_result164[23]^and_result164[24]^and_result164[25]^and_result164[26]^and_result164[27]^and_result164[28]^and_result164[29]^and_result164[30]^and_result164[31]^and_result164[32]^and_result164[33]^and_result164[34]^and_result164[35]^and_result164[36]^and_result164[37]^and_result164[38]^and_result164[39]^and_result164[40]^and_result164[41]^and_result164[42]^and_result164[43]^and_result164[44]^and_result164[45]^and_result164[46]^and_result164[47]^and_result164[48]^and_result164[49]^and_result164[50]^and_result164[51]^and_result164[52]^and_result164[53]^and_result164[54]^and_result164[55]^and_result164[56]^and_result164[57]^and_result164[58]^and_result164[59]^and_result164[60]^and_result164[61]^and_result164[62]^and_result164[63]^and_result164[64]^and_result164[65]^and_result164[66]^and_result164[67]^and_result164[68]^and_result164[69]^and_result164[70]^and_result164[71]^and_result164[72]^and_result164[73]^and_result164[74]^and_result164[75]^and_result164[76]^and_result164[77]^and_result164[78]^and_result164[79]^and_result164[80]^and_result164[81]^and_result164[82]^and_result164[83]^and_result164[84]^and_result164[85]^and_result164[86]^and_result164[87]^and_result164[88]^and_result164[89]^and_result164[90]^and_result164[91]^and_result164[92]^and_result164[93]^and_result164[94]^and_result164[95]^and_result164[96]^and_result164[97]^and_result164[98]^and_result164[99]^and_result164[100]^and_result164[101]^and_result164[102]^and_result164[103]^and_result164[104]^and_result164[105]^and_result164[106]^and_result164[107]^and_result164[108]^and_result164[109]^and_result164[110]^and_result164[111]^and_result164[112]^and_result164[113]^and_result164[114]^and_result164[115]^and_result164[116]^and_result164[117]^and_result164[118]^and_result164[119]^and_result164[120]^and_result164[121]^and_result164[122]^and_result164[123]^and_result164[124]^and_result164[125]^and_result164[126]^and_result164[127]^and_result164[128]^and_result164[129]^and_result164[130]^and_result164[131]^and_result164[132]^and_result164[133]^and_result164[134]^and_result164[135]^and_result164[136]^and_result164[137]^and_result164[138]^and_result164[139]^and_result164[140]^and_result164[141]^and_result164[142]^and_result164[143]^and_result164[144]^and_result164[145]^and_result164[146]^and_result164[147]^and_result164[148]^and_result164[149]^and_result164[150]^and_result164[151]^and_result164[152]^and_result164[153]^and_result164[154]^and_result164[155]^and_result164[156]^and_result164[157]^and_result164[158]^and_result164[159]^and_result164[160]^and_result164[161]^and_result164[162]^and_result164[163]^and_result164[164]^and_result164[165]^and_result164[166]^and_result164[167]^and_result164[168]^and_result164[169]^and_result164[170]^and_result164[171]^and_result164[172]^and_result164[173]^and_result164[174]^and_result164[175]^and_result164[176]^and_result164[177]^and_result164[178]^and_result164[179]^and_result164[180]^and_result164[181]^and_result164[182]^and_result164[183]^and_result164[184]^and_result164[185]^and_result164[186]^and_result164[187]^and_result164[188]^and_result164[189]^and_result164[190]^and_result164[191]^and_result164[192]^and_result164[193]^and_result164[194]^and_result164[195]^and_result164[196]^and_result164[197]^and_result164[198]^and_result164[199]^and_result164[200]^and_result164[201]^and_result164[202]^and_result164[203]^and_result164[204]^and_result164[205]^and_result164[206]^and_result164[207]^and_result164[208]^and_result164[209]^and_result164[210]^and_result164[211]^and_result164[212]^and_result164[213]^and_result164[214]^and_result164[215]^and_result164[216]^and_result164[217]^and_result164[218]^and_result164[219]^and_result164[220]^and_result164[221]^and_result164[222]^and_result164[223]^and_result164[224]^and_result164[225]^and_result164[226]^and_result164[227]^and_result164[228]^and_result164[229]^and_result164[230]^and_result164[231]^and_result164[232]^and_result164[233]^and_result164[234]^and_result164[235]^and_result164[236]^and_result164[237]^and_result164[238]^and_result164[239]^and_result164[240]^and_result164[241]^and_result164[242]^and_result164[243]^and_result164[244]^and_result164[245]^and_result164[246]^and_result164[247]^and_result164[248]^and_result164[249]^and_result164[250]^and_result164[251]^and_result164[252]^and_result164[253]^and_result164[254];
assign key[165]=and_result165[0]^and_result165[1]^and_result165[2]^and_result165[3]^and_result165[4]^and_result165[5]^and_result165[6]^and_result165[7]^and_result165[8]^and_result165[9]^and_result165[10]^and_result165[11]^and_result165[12]^and_result165[13]^and_result165[14]^and_result165[15]^and_result165[16]^and_result165[17]^and_result165[18]^and_result165[19]^and_result165[20]^and_result165[21]^and_result165[22]^and_result165[23]^and_result165[24]^and_result165[25]^and_result165[26]^and_result165[27]^and_result165[28]^and_result165[29]^and_result165[30]^and_result165[31]^and_result165[32]^and_result165[33]^and_result165[34]^and_result165[35]^and_result165[36]^and_result165[37]^and_result165[38]^and_result165[39]^and_result165[40]^and_result165[41]^and_result165[42]^and_result165[43]^and_result165[44]^and_result165[45]^and_result165[46]^and_result165[47]^and_result165[48]^and_result165[49]^and_result165[50]^and_result165[51]^and_result165[52]^and_result165[53]^and_result165[54]^and_result165[55]^and_result165[56]^and_result165[57]^and_result165[58]^and_result165[59]^and_result165[60]^and_result165[61]^and_result165[62]^and_result165[63]^and_result165[64]^and_result165[65]^and_result165[66]^and_result165[67]^and_result165[68]^and_result165[69]^and_result165[70]^and_result165[71]^and_result165[72]^and_result165[73]^and_result165[74]^and_result165[75]^and_result165[76]^and_result165[77]^and_result165[78]^and_result165[79]^and_result165[80]^and_result165[81]^and_result165[82]^and_result165[83]^and_result165[84]^and_result165[85]^and_result165[86]^and_result165[87]^and_result165[88]^and_result165[89]^and_result165[90]^and_result165[91]^and_result165[92]^and_result165[93]^and_result165[94]^and_result165[95]^and_result165[96]^and_result165[97]^and_result165[98]^and_result165[99]^and_result165[100]^and_result165[101]^and_result165[102]^and_result165[103]^and_result165[104]^and_result165[105]^and_result165[106]^and_result165[107]^and_result165[108]^and_result165[109]^and_result165[110]^and_result165[111]^and_result165[112]^and_result165[113]^and_result165[114]^and_result165[115]^and_result165[116]^and_result165[117]^and_result165[118]^and_result165[119]^and_result165[120]^and_result165[121]^and_result165[122]^and_result165[123]^and_result165[124]^and_result165[125]^and_result165[126]^and_result165[127]^and_result165[128]^and_result165[129]^and_result165[130]^and_result165[131]^and_result165[132]^and_result165[133]^and_result165[134]^and_result165[135]^and_result165[136]^and_result165[137]^and_result165[138]^and_result165[139]^and_result165[140]^and_result165[141]^and_result165[142]^and_result165[143]^and_result165[144]^and_result165[145]^and_result165[146]^and_result165[147]^and_result165[148]^and_result165[149]^and_result165[150]^and_result165[151]^and_result165[152]^and_result165[153]^and_result165[154]^and_result165[155]^and_result165[156]^and_result165[157]^and_result165[158]^and_result165[159]^and_result165[160]^and_result165[161]^and_result165[162]^and_result165[163]^and_result165[164]^and_result165[165]^and_result165[166]^and_result165[167]^and_result165[168]^and_result165[169]^and_result165[170]^and_result165[171]^and_result165[172]^and_result165[173]^and_result165[174]^and_result165[175]^and_result165[176]^and_result165[177]^and_result165[178]^and_result165[179]^and_result165[180]^and_result165[181]^and_result165[182]^and_result165[183]^and_result165[184]^and_result165[185]^and_result165[186]^and_result165[187]^and_result165[188]^and_result165[189]^and_result165[190]^and_result165[191]^and_result165[192]^and_result165[193]^and_result165[194]^and_result165[195]^and_result165[196]^and_result165[197]^and_result165[198]^and_result165[199]^and_result165[200]^and_result165[201]^and_result165[202]^and_result165[203]^and_result165[204]^and_result165[205]^and_result165[206]^and_result165[207]^and_result165[208]^and_result165[209]^and_result165[210]^and_result165[211]^and_result165[212]^and_result165[213]^and_result165[214]^and_result165[215]^and_result165[216]^and_result165[217]^and_result165[218]^and_result165[219]^and_result165[220]^and_result165[221]^and_result165[222]^and_result165[223]^and_result165[224]^and_result165[225]^and_result165[226]^and_result165[227]^and_result165[228]^and_result165[229]^and_result165[230]^and_result165[231]^and_result165[232]^and_result165[233]^and_result165[234]^and_result165[235]^and_result165[236]^and_result165[237]^and_result165[238]^and_result165[239]^and_result165[240]^and_result165[241]^and_result165[242]^and_result165[243]^and_result165[244]^and_result165[245]^and_result165[246]^and_result165[247]^and_result165[248]^and_result165[249]^and_result165[250]^and_result165[251]^and_result165[252]^and_result165[253]^and_result165[254];
assign key[166]=and_result166[0]^and_result166[1]^and_result166[2]^and_result166[3]^and_result166[4]^and_result166[5]^and_result166[6]^and_result166[7]^and_result166[8]^and_result166[9]^and_result166[10]^and_result166[11]^and_result166[12]^and_result166[13]^and_result166[14]^and_result166[15]^and_result166[16]^and_result166[17]^and_result166[18]^and_result166[19]^and_result166[20]^and_result166[21]^and_result166[22]^and_result166[23]^and_result166[24]^and_result166[25]^and_result166[26]^and_result166[27]^and_result166[28]^and_result166[29]^and_result166[30]^and_result166[31]^and_result166[32]^and_result166[33]^and_result166[34]^and_result166[35]^and_result166[36]^and_result166[37]^and_result166[38]^and_result166[39]^and_result166[40]^and_result166[41]^and_result166[42]^and_result166[43]^and_result166[44]^and_result166[45]^and_result166[46]^and_result166[47]^and_result166[48]^and_result166[49]^and_result166[50]^and_result166[51]^and_result166[52]^and_result166[53]^and_result166[54]^and_result166[55]^and_result166[56]^and_result166[57]^and_result166[58]^and_result166[59]^and_result166[60]^and_result166[61]^and_result166[62]^and_result166[63]^and_result166[64]^and_result166[65]^and_result166[66]^and_result166[67]^and_result166[68]^and_result166[69]^and_result166[70]^and_result166[71]^and_result166[72]^and_result166[73]^and_result166[74]^and_result166[75]^and_result166[76]^and_result166[77]^and_result166[78]^and_result166[79]^and_result166[80]^and_result166[81]^and_result166[82]^and_result166[83]^and_result166[84]^and_result166[85]^and_result166[86]^and_result166[87]^and_result166[88]^and_result166[89]^and_result166[90]^and_result166[91]^and_result166[92]^and_result166[93]^and_result166[94]^and_result166[95]^and_result166[96]^and_result166[97]^and_result166[98]^and_result166[99]^and_result166[100]^and_result166[101]^and_result166[102]^and_result166[103]^and_result166[104]^and_result166[105]^and_result166[106]^and_result166[107]^and_result166[108]^and_result166[109]^and_result166[110]^and_result166[111]^and_result166[112]^and_result166[113]^and_result166[114]^and_result166[115]^and_result166[116]^and_result166[117]^and_result166[118]^and_result166[119]^and_result166[120]^and_result166[121]^and_result166[122]^and_result166[123]^and_result166[124]^and_result166[125]^and_result166[126]^and_result166[127]^and_result166[128]^and_result166[129]^and_result166[130]^and_result166[131]^and_result166[132]^and_result166[133]^and_result166[134]^and_result166[135]^and_result166[136]^and_result166[137]^and_result166[138]^and_result166[139]^and_result166[140]^and_result166[141]^and_result166[142]^and_result166[143]^and_result166[144]^and_result166[145]^and_result166[146]^and_result166[147]^and_result166[148]^and_result166[149]^and_result166[150]^and_result166[151]^and_result166[152]^and_result166[153]^and_result166[154]^and_result166[155]^and_result166[156]^and_result166[157]^and_result166[158]^and_result166[159]^and_result166[160]^and_result166[161]^and_result166[162]^and_result166[163]^and_result166[164]^and_result166[165]^and_result166[166]^and_result166[167]^and_result166[168]^and_result166[169]^and_result166[170]^and_result166[171]^and_result166[172]^and_result166[173]^and_result166[174]^and_result166[175]^and_result166[176]^and_result166[177]^and_result166[178]^and_result166[179]^and_result166[180]^and_result166[181]^and_result166[182]^and_result166[183]^and_result166[184]^and_result166[185]^and_result166[186]^and_result166[187]^and_result166[188]^and_result166[189]^and_result166[190]^and_result166[191]^and_result166[192]^and_result166[193]^and_result166[194]^and_result166[195]^and_result166[196]^and_result166[197]^and_result166[198]^and_result166[199]^and_result166[200]^and_result166[201]^and_result166[202]^and_result166[203]^and_result166[204]^and_result166[205]^and_result166[206]^and_result166[207]^and_result166[208]^and_result166[209]^and_result166[210]^and_result166[211]^and_result166[212]^and_result166[213]^and_result166[214]^and_result166[215]^and_result166[216]^and_result166[217]^and_result166[218]^and_result166[219]^and_result166[220]^and_result166[221]^and_result166[222]^and_result166[223]^and_result166[224]^and_result166[225]^and_result166[226]^and_result166[227]^and_result166[228]^and_result166[229]^and_result166[230]^and_result166[231]^and_result166[232]^and_result166[233]^and_result166[234]^and_result166[235]^and_result166[236]^and_result166[237]^and_result166[238]^and_result166[239]^and_result166[240]^and_result166[241]^and_result166[242]^and_result166[243]^and_result166[244]^and_result166[245]^and_result166[246]^and_result166[247]^and_result166[248]^and_result166[249]^and_result166[250]^and_result166[251]^and_result166[252]^and_result166[253]^and_result166[254];
assign key[167]=and_result167[0]^and_result167[1]^and_result167[2]^and_result167[3]^and_result167[4]^and_result167[5]^and_result167[6]^and_result167[7]^and_result167[8]^and_result167[9]^and_result167[10]^and_result167[11]^and_result167[12]^and_result167[13]^and_result167[14]^and_result167[15]^and_result167[16]^and_result167[17]^and_result167[18]^and_result167[19]^and_result167[20]^and_result167[21]^and_result167[22]^and_result167[23]^and_result167[24]^and_result167[25]^and_result167[26]^and_result167[27]^and_result167[28]^and_result167[29]^and_result167[30]^and_result167[31]^and_result167[32]^and_result167[33]^and_result167[34]^and_result167[35]^and_result167[36]^and_result167[37]^and_result167[38]^and_result167[39]^and_result167[40]^and_result167[41]^and_result167[42]^and_result167[43]^and_result167[44]^and_result167[45]^and_result167[46]^and_result167[47]^and_result167[48]^and_result167[49]^and_result167[50]^and_result167[51]^and_result167[52]^and_result167[53]^and_result167[54]^and_result167[55]^and_result167[56]^and_result167[57]^and_result167[58]^and_result167[59]^and_result167[60]^and_result167[61]^and_result167[62]^and_result167[63]^and_result167[64]^and_result167[65]^and_result167[66]^and_result167[67]^and_result167[68]^and_result167[69]^and_result167[70]^and_result167[71]^and_result167[72]^and_result167[73]^and_result167[74]^and_result167[75]^and_result167[76]^and_result167[77]^and_result167[78]^and_result167[79]^and_result167[80]^and_result167[81]^and_result167[82]^and_result167[83]^and_result167[84]^and_result167[85]^and_result167[86]^and_result167[87]^and_result167[88]^and_result167[89]^and_result167[90]^and_result167[91]^and_result167[92]^and_result167[93]^and_result167[94]^and_result167[95]^and_result167[96]^and_result167[97]^and_result167[98]^and_result167[99]^and_result167[100]^and_result167[101]^and_result167[102]^and_result167[103]^and_result167[104]^and_result167[105]^and_result167[106]^and_result167[107]^and_result167[108]^and_result167[109]^and_result167[110]^and_result167[111]^and_result167[112]^and_result167[113]^and_result167[114]^and_result167[115]^and_result167[116]^and_result167[117]^and_result167[118]^and_result167[119]^and_result167[120]^and_result167[121]^and_result167[122]^and_result167[123]^and_result167[124]^and_result167[125]^and_result167[126]^and_result167[127]^and_result167[128]^and_result167[129]^and_result167[130]^and_result167[131]^and_result167[132]^and_result167[133]^and_result167[134]^and_result167[135]^and_result167[136]^and_result167[137]^and_result167[138]^and_result167[139]^and_result167[140]^and_result167[141]^and_result167[142]^and_result167[143]^and_result167[144]^and_result167[145]^and_result167[146]^and_result167[147]^and_result167[148]^and_result167[149]^and_result167[150]^and_result167[151]^and_result167[152]^and_result167[153]^and_result167[154]^and_result167[155]^and_result167[156]^and_result167[157]^and_result167[158]^and_result167[159]^and_result167[160]^and_result167[161]^and_result167[162]^and_result167[163]^and_result167[164]^and_result167[165]^and_result167[166]^and_result167[167]^and_result167[168]^and_result167[169]^and_result167[170]^and_result167[171]^and_result167[172]^and_result167[173]^and_result167[174]^and_result167[175]^and_result167[176]^and_result167[177]^and_result167[178]^and_result167[179]^and_result167[180]^and_result167[181]^and_result167[182]^and_result167[183]^and_result167[184]^and_result167[185]^and_result167[186]^and_result167[187]^and_result167[188]^and_result167[189]^and_result167[190]^and_result167[191]^and_result167[192]^and_result167[193]^and_result167[194]^and_result167[195]^and_result167[196]^and_result167[197]^and_result167[198]^and_result167[199]^and_result167[200]^and_result167[201]^and_result167[202]^and_result167[203]^and_result167[204]^and_result167[205]^and_result167[206]^and_result167[207]^and_result167[208]^and_result167[209]^and_result167[210]^and_result167[211]^and_result167[212]^and_result167[213]^and_result167[214]^and_result167[215]^and_result167[216]^and_result167[217]^and_result167[218]^and_result167[219]^and_result167[220]^and_result167[221]^and_result167[222]^and_result167[223]^and_result167[224]^and_result167[225]^and_result167[226]^and_result167[227]^and_result167[228]^and_result167[229]^and_result167[230]^and_result167[231]^and_result167[232]^and_result167[233]^and_result167[234]^and_result167[235]^and_result167[236]^and_result167[237]^and_result167[238]^and_result167[239]^and_result167[240]^and_result167[241]^and_result167[242]^and_result167[243]^and_result167[244]^and_result167[245]^and_result167[246]^and_result167[247]^and_result167[248]^and_result167[249]^and_result167[250]^and_result167[251]^and_result167[252]^and_result167[253]^and_result167[254];
assign key[168]=and_result168[0]^and_result168[1]^and_result168[2]^and_result168[3]^and_result168[4]^and_result168[5]^and_result168[6]^and_result168[7]^and_result168[8]^and_result168[9]^and_result168[10]^and_result168[11]^and_result168[12]^and_result168[13]^and_result168[14]^and_result168[15]^and_result168[16]^and_result168[17]^and_result168[18]^and_result168[19]^and_result168[20]^and_result168[21]^and_result168[22]^and_result168[23]^and_result168[24]^and_result168[25]^and_result168[26]^and_result168[27]^and_result168[28]^and_result168[29]^and_result168[30]^and_result168[31]^and_result168[32]^and_result168[33]^and_result168[34]^and_result168[35]^and_result168[36]^and_result168[37]^and_result168[38]^and_result168[39]^and_result168[40]^and_result168[41]^and_result168[42]^and_result168[43]^and_result168[44]^and_result168[45]^and_result168[46]^and_result168[47]^and_result168[48]^and_result168[49]^and_result168[50]^and_result168[51]^and_result168[52]^and_result168[53]^and_result168[54]^and_result168[55]^and_result168[56]^and_result168[57]^and_result168[58]^and_result168[59]^and_result168[60]^and_result168[61]^and_result168[62]^and_result168[63]^and_result168[64]^and_result168[65]^and_result168[66]^and_result168[67]^and_result168[68]^and_result168[69]^and_result168[70]^and_result168[71]^and_result168[72]^and_result168[73]^and_result168[74]^and_result168[75]^and_result168[76]^and_result168[77]^and_result168[78]^and_result168[79]^and_result168[80]^and_result168[81]^and_result168[82]^and_result168[83]^and_result168[84]^and_result168[85]^and_result168[86]^and_result168[87]^and_result168[88]^and_result168[89]^and_result168[90]^and_result168[91]^and_result168[92]^and_result168[93]^and_result168[94]^and_result168[95]^and_result168[96]^and_result168[97]^and_result168[98]^and_result168[99]^and_result168[100]^and_result168[101]^and_result168[102]^and_result168[103]^and_result168[104]^and_result168[105]^and_result168[106]^and_result168[107]^and_result168[108]^and_result168[109]^and_result168[110]^and_result168[111]^and_result168[112]^and_result168[113]^and_result168[114]^and_result168[115]^and_result168[116]^and_result168[117]^and_result168[118]^and_result168[119]^and_result168[120]^and_result168[121]^and_result168[122]^and_result168[123]^and_result168[124]^and_result168[125]^and_result168[126]^and_result168[127]^and_result168[128]^and_result168[129]^and_result168[130]^and_result168[131]^and_result168[132]^and_result168[133]^and_result168[134]^and_result168[135]^and_result168[136]^and_result168[137]^and_result168[138]^and_result168[139]^and_result168[140]^and_result168[141]^and_result168[142]^and_result168[143]^and_result168[144]^and_result168[145]^and_result168[146]^and_result168[147]^and_result168[148]^and_result168[149]^and_result168[150]^and_result168[151]^and_result168[152]^and_result168[153]^and_result168[154]^and_result168[155]^and_result168[156]^and_result168[157]^and_result168[158]^and_result168[159]^and_result168[160]^and_result168[161]^and_result168[162]^and_result168[163]^and_result168[164]^and_result168[165]^and_result168[166]^and_result168[167]^and_result168[168]^and_result168[169]^and_result168[170]^and_result168[171]^and_result168[172]^and_result168[173]^and_result168[174]^and_result168[175]^and_result168[176]^and_result168[177]^and_result168[178]^and_result168[179]^and_result168[180]^and_result168[181]^and_result168[182]^and_result168[183]^and_result168[184]^and_result168[185]^and_result168[186]^and_result168[187]^and_result168[188]^and_result168[189]^and_result168[190]^and_result168[191]^and_result168[192]^and_result168[193]^and_result168[194]^and_result168[195]^and_result168[196]^and_result168[197]^and_result168[198]^and_result168[199]^and_result168[200]^and_result168[201]^and_result168[202]^and_result168[203]^and_result168[204]^and_result168[205]^and_result168[206]^and_result168[207]^and_result168[208]^and_result168[209]^and_result168[210]^and_result168[211]^and_result168[212]^and_result168[213]^and_result168[214]^and_result168[215]^and_result168[216]^and_result168[217]^and_result168[218]^and_result168[219]^and_result168[220]^and_result168[221]^and_result168[222]^and_result168[223]^and_result168[224]^and_result168[225]^and_result168[226]^and_result168[227]^and_result168[228]^and_result168[229]^and_result168[230]^and_result168[231]^and_result168[232]^and_result168[233]^and_result168[234]^and_result168[235]^and_result168[236]^and_result168[237]^and_result168[238]^and_result168[239]^and_result168[240]^and_result168[241]^and_result168[242]^and_result168[243]^and_result168[244]^and_result168[245]^and_result168[246]^and_result168[247]^and_result168[248]^and_result168[249]^and_result168[250]^and_result168[251]^and_result168[252]^and_result168[253]^and_result168[254];
assign key[169]=and_result169[0]^and_result169[1]^and_result169[2]^and_result169[3]^and_result169[4]^and_result169[5]^and_result169[6]^and_result169[7]^and_result169[8]^and_result169[9]^and_result169[10]^and_result169[11]^and_result169[12]^and_result169[13]^and_result169[14]^and_result169[15]^and_result169[16]^and_result169[17]^and_result169[18]^and_result169[19]^and_result169[20]^and_result169[21]^and_result169[22]^and_result169[23]^and_result169[24]^and_result169[25]^and_result169[26]^and_result169[27]^and_result169[28]^and_result169[29]^and_result169[30]^and_result169[31]^and_result169[32]^and_result169[33]^and_result169[34]^and_result169[35]^and_result169[36]^and_result169[37]^and_result169[38]^and_result169[39]^and_result169[40]^and_result169[41]^and_result169[42]^and_result169[43]^and_result169[44]^and_result169[45]^and_result169[46]^and_result169[47]^and_result169[48]^and_result169[49]^and_result169[50]^and_result169[51]^and_result169[52]^and_result169[53]^and_result169[54]^and_result169[55]^and_result169[56]^and_result169[57]^and_result169[58]^and_result169[59]^and_result169[60]^and_result169[61]^and_result169[62]^and_result169[63]^and_result169[64]^and_result169[65]^and_result169[66]^and_result169[67]^and_result169[68]^and_result169[69]^and_result169[70]^and_result169[71]^and_result169[72]^and_result169[73]^and_result169[74]^and_result169[75]^and_result169[76]^and_result169[77]^and_result169[78]^and_result169[79]^and_result169[80]^and_result169[81]^and_result169[82]^and_result169[83]^and_result169[84]^and_result169[85]^and_result169[86]^and_result169[87]^and_result169[88]^and_result169[89]^and_result169[90]^and_result169[91]^and_result169[92]^and_result169[93]^and_result169[94]^and_result169[95]^and_result169[96]^and_result169[97]^and_result169[98]^and_result169[99]^and_result169[100]^and_result169[101]^and_result169[102]^and_result169[103]^and_result169[104]^and_result169[105]^and_result169[106]^and_result169[107]^and_result169[108]^and_result169[109]^and_result169[110]^and_result169[111]^and_result169[112]^and_result169[113]^and_result169[114]^and_result169[115]^and_result169[116]^and_result169[117]^and_result169[118]^and_result169[119]^and_result169[120]^and_result169[121]^and_result169[122]^and_result169[123]^and_result169[124]^and_result169[125]^and_result169[126]^and_result169[127]^and_result169[128]^and_result169[129]^and_result169[130]^and_result169[131]^and_result169[132]^and_result169[133]^and_result169[134]^and_result169[135]^and_result169[136]^and_result169[137]^and_result169[138]^and_result169[139]^and_result169[140]^and_result169[141]^and_result169[142]^and_result169[143]^and_result169[144]^and_result169[145]^and_result169[146]^and_result169[147]^and_result169[148]^and_result169[149]^and_result169[150]^and_result169[151]^and_result169[152]^and_result169[153]^and_result169[154]^and_result169[155]^and_result169[156]^and_result169[157]^and_result169[158]^and_result169[159]^and_result169[160]^and_result169[161]^and_result169[162]^and_result169[163]^and_result169[164]^and_result169[165]^and_result169[166]^and_result169[167]^and_result169[168]^and_result169[169]^and_result169[170]^and_result169[171]^and_result169[172]^and_result169[173]^and_result169[174]^and_result169[175]^and_result169[176]^and_result169[177]^and_result169[178]^and_result169[179]^and_result169[180]^and_result169[181]^and_result169[182]^and_result169[183]^and_result169[184]^and_result169[185]^and_result169[186]^and_result169[187]^and_result169[188]^and_result169[189]^and_result169[190]^and_result169[191]^and_result169[192]^and_result169[193]^and_result169[194]^and_result169[195]^and_result169[196]^and_result169[197]^and_result169[198]^and_result169[199]^and_result169[200]^and_result169[201]^and_result169[202]^and_result169[203]^and_result169[204]^and_result169[205]^and_result169[206]^and_result169[207]^and_result169[208]^and_result169[209]^and_result169[210]^and_result169[211]^and_result169[212]^and_result169[213]^and_result169[214]^and_result169[215]^and_result169[216]^and_result169[217]^and_result169[218]^and_result169[219]^and_result169[220]^and_result169[221]^and_result169[222]^and_result169[223]^and_result169[224]^and_result169[225]^and_result169[226]^and_result169[227]^and_result169[228]^and_result169[229]^and_result169[230]^and_result169[231]^and_result169[232]^and_result169[233]^and_result169[234]^and_result169[235]^and_result169[236]^and_result169[237]^and_result169[238]^and_result169[239]^and_result169[240]^and_result169[241]^and_result169[242]^and_result169[243]^and_result169[244]^and_result169[245]^and_result169[246]^and_result169[247]^and_result169[248]^and_result169[249]^and_result169[250]^and_result169[251]^and_result169[252]^and_result169[253]^and_result169[254];
assign key[170]=and_result170[0]^and_result170[1]^and_result170[2]^and_result170[3]^and_result170[4]^and_result170[5]^and_result170[6]^and_result170[7]^and_result170[8]^and_result170[9]^and_result170[10]^and_result170[11]^and_result170[12]^and_result170[13]^and_result170[14]^and_result170[15]^and_result170[16]^and_result170[17]^and_result170[18]^and_result170[19]^and_result170[20]^and_result170[21]^and_result170[22]^and_result170[23]^and_result170[24]^and_result170[25]^and_result170[26]^and_result170[27]^and_result170[28]^and_result170[29]^and_result170[30]^and_result170[31]^and_result170[32]^and_result170[33]^and_result170[34]^and_result170[35]^and_result170[36]^and_result170[37]^and_result170[38]^and_result170[39]^and_result170[40]^and_result170[41]^and_result170[42]^and_result170[43]^and_result170[44]^and_result170[45]^and_result170[46]^and_result170[47]^and_result170[48]^and_result170[49]^and_result170[50]^and_result170[51]^and_result170[52]^and_result170[53]^and_result170[54]^and_result170[55]^and_result170[56]^and_result170[57]^and_result170[58]^and_result170[59]^and_result170[60]^and_result170[61]^and_result170[62]^and_result170[63]^and_result170[64]^and_result170[65]^and_result170[66]^and_result170[67]^and_result170[68]^and_result170[69]^and_result170[70]^and_result170[71]^and_result170[72]^and_result170[73]^and_result170[74]^and_result170[75]^and_result170[76]^and_result170[77]^and_result170[78]^and_result170[79]^and_result170[80]^and_result170[81]^and_result170[82]^and_result170[83]^and_result170[84]^and_result170[85]^and_result170[86]^and_result170[87]^and_result170[88]^and_result170[89]^and_result170[90]^and_result170[91]^and_result170[92]^and_result170[93]^and_result170[94]^and_result170[95]^and_result170[96]^and_result170[97]^and_result170[98]^and_result170[99]^and_result170[100]^and_result170[101]^and_result170[102]^and_result170[103]^and_result170[104]^and_result170[105]^and_result170[106]^and_result170[107]^and_result170[108]^and_result170[109]^and_result170[110]^and_result170[111]^and_result170[112]^and_result170[113]^and_result170[114]^and_result170[115]^and_result170[116]^and_result170[117]^and_result170[118]^and_result170[119]^and_result170[120]^and_result170[121]^and_result170[122]^and_result170[123]^and_result170[124]^and_result170[125]^and_result170[126]^and_result170[127]^and_result170[128]^and_result170[129]^and_result170[130]^and_result170[131]^and_result170[132]^and_result170[133]^and_result170[134]^and_result170[135]^and_result170[136]^and_result170[137]^and_result170[138]^and_result170[139]^and_result170[140]^and_result170[141]^and_result170[142]^and_result170[143]^and_result170[144]^and_result170[145]^and_result170[146]^and_result170[147]^and_result170[148]^and_result170[149]^and_result170[150]^and_result170[151]^and_result170[152]^and_result170[153]^and_result170[154]^and_result170[155]^and_result170[156]^and_result170[157]^and_result170[158]^and_result170[159]^and_result170[160]^and_result170[161]^and_result170[162]^and_result170[163]^and_result170[164]^and_result170[165]^and_result170[166]^and_result170[167]^and_result170[168]^and_result170[169]^and_result170[170]^and_result170[171]^and_result170[172]^and_result170[173]^and_result170[174]^and_result170[175]^and_result170[176]^and_result170[177]^and_result170[178]^and_result170[179]^and_result170[180]^and_result170[181]^and_result170[182]^and_result170[183]^and_result170[184]^and_result170[185]^and_result170[186]^and_result170[187]^and_result170[188]^and_result170[189]^and_result170[190]^and_result170[191]^and_result170[192]^and_result170[193]^and_result170[194]^and_result170[195]^and_result170[196]^and_result170[197]^and_result170[198]^and_result170[199]^and_result170[200]^and_result170[201]^and_result170[202]^and_result170[203]^and_result170[204]^and_result170[205]^and_result170[206]^and_result170[207]^and_result170[208]^and_result170[209]^and_result170[210]^and_result170[211]^and_result170[212]^and_result170[213]^and_result170[214]^and_result170[215]^and_result170[216]^and_result170[217]^and_result170[218]^and_result170[219]^and_result170[220]^and_result170[221]^and_result170[222]^and_result170[223]^and_result170[224]^and_result170[225]^and_result170[226]^and_result170[227]^and_result170[228]^and_result170[229]^and_result170[230]^and_result170[231]^and_result170[232]^and_result170[233]^and_result170[234]^and_result170[235]^and_result170[236]^and_result170[237]^and_result170[238]^and_result170[239]^and_result170[240]^and_result170[241]^and_result170[242]^and_result170[243]^and_result170[244]^and_result170[245]^and_result170[246]^and_result170[247]^and_result170[248]^and_result170[249]^and_result170[250]^and_result170[251]^and_result170[252]^and_result170[253]^and_result170[254];
assign key[171]=and_result171[0]^and_result171[1]^and_result171[2]^and_result171[3]^and_result171[4]^and_result171[5]^and_result171[6]^and_result171[7]^and_result171[8]^and_result171[9]^and_result171[10]^and_result171[11]^and_result171[12]^and_result171[13]^and_result171[14]^and_result171[15]^and_result171[16]^and_result171[17]^and_result171[18]^and_result171[19]^and_result171[20]^and_result171[21]^and_result171[22]^and_result171[23]^and_result171[24]^and_result171[25]^and_result171[26]^and_result171[27]^and_result171[28]^and_result171[29]^and_result171[30]^and_result171[31]^and_result171[32]^and_result171[33]^and_result171[34]^and_result171[35]^and_result171[36]^and_result171[37]^and_result171[38]^and_result171[39]^and_result171[40]^and_result171[41]^and_result171[42]^and_result171[43]^and_result171[44]^and_result171[45]^and_result171[46]^and_result171[47]^and_result171[48]^and_result171[49]^and_result171[50]^and_result171[51]^and_result171[52]^and_result171[53]^and_result171[54]^and_result171[55]^and_result171[56]^and_result171[57]^and_result171[58]^and_result171[59]^and_result171[60]^and_result171[61]^and_result171[62]^and_result171[63]^and_result171[64]^and_result171[65]^and_result171[66]^and_result171[67]^and_result171[68]^and_result171[69]^and_result171[70]^and_result171[71]^and_result171[72]^and_result171[73]^and_result171[74]^and_result171[75]^and_result171[76]^and_result171[77]^and_result171[78]^and_result171[79]^and_result171[80]^and_result171[81]^and_result171[82]^and_result171[83]^and_result171[84]^and_result171[85]^and_result171[86]^and_result171[87]^and_result171[88]^and_result171[89]^and_result171[90]^and_result171[91]^and_result171[92]^and_result171[93]^and_result171[94]^and_result171[95]^and_result171[96]^and_result171[97]^and_result171[98]^and_result171[99]^and_result171[100]^and_result171[101]^and_result171[102]^and_result171[103]^and_result171[104]^and_result171[105]^and_result171[106]^and_result171[107]^and_result171[108]^and_result171[109]^and_result171[110]^and_result171[111]^and_result171[112]^and_result171[113]^and_result171[114]^and_result171[115]^and_result171[116]^and_result171[117]^and_result171[118]^and_result171[119]^and_result171[120]^and_result171[121]^and_result171[122]^and_result171[123]^and_result171[124]^and_result171[125]^and_result171[126]^and_result171[127]^and_result171[128]^and_result171[129]^and_result171[130]^and_result171[131]^and_result171[132]^and_result171[133]^and_result171[134]^and_result171[135]^and_result171[136]^and_result171[137]^and_result171[138]^and_result171[139]^and_result171[140]^and_result171[141]^and_result171[142]^and_result171[143]^and_result171[144]^and_result171[145]^and_result171[146]^and_result171[147]^and_result171[148]^and_result171[149]^and_result171[150]^and_result171[151]^and_result171[152]^and_result171[153]^and_result171[154]^and_result171[155]^and_result171[156]^and_result171[157]^and_result171[158]^and_result171[159]^and_result171[160]^and_result171[161]^and_result171[162]^and_result171[163]^and_result171[164]^and_result171[165]^and_result171[166]^and_result171[167]^and_result171[168]^and_result171[169]^and_result171[170]^and_result171[171]^and_result171[172]^and_result171[173]^and_result171[174]^and_result171[175]^and_result171[176]^and_result171[177]^and_result171[178]^and_result171[179]^and_result171[180]^and_result171[181]^and_result171[182]^and_result171[183]^and_result171[184]^and_result171[185]^and_result171[186]^and_result171[187]^and_result171[188]^and_result171[189]^and_result171[190]^and_result171[191]^and_result171[192]^and_result171[193]^and_result171[194]^and_result171[195]^and_result171[196]^and_result171[197]^and_result171[198]^and_result171[199]^and_result171[200]^and_result171[201]^and_result171[202]^and_result171[203]^and_result171[204]^and_result171[205]^and_result171[206]^and_result171[207]^and_result171[208]^and_result171[209]^and_result171[210]^and_result171[211]^and_result171[212]^and_result171[213]^and_result171[214]^and_result171[215]^and_result171[216]^and_result171[217]^and_result171[218]^and_result171[219]^and_result171[220]^and_result171[221]^and_result171[222]^and_result171[223]^and_result171[224]^and_result171[225]^and_result171[226]^and_result171[227]^and_result171[228]^and_result171[229]^and_result171[230]^and_result171[231]^and_result171[232]^and_result171[233]^and_result171[234]^and_result171[235]^and_result171[236]^and_result171[237]^and_result171[238]^and_result171[239]^and_result171[240]^and_result171[241]^and_result171[242]^and_result171[243]^and_result171[244]^and_result171[245]^and_result171[246]^and_result171[247]^and_result171[248]^and_result171[249]^and_result171[250]^and_result171[251]^and_result171[252]^and_result171[253]^and_result171[254];
assign key[172]=and_result172[0]^and_result172[1]^and_result172[2]^and_result172[3]^and_result172[4]^and_result172[5]^and_result172[6]^and_result172[7]^and_result172[8]^and_result172[9]^and_result172[10]^and_result172[11]^and_result172[12]^and_result172[13]^and_result172[14]^and_result172[15]^and_result172[16]^and_result172[17]^and_result172[18]^and_result172[19]^and_result172[20]^and_result172[21]^and_result172[22]^and_result172[23]^and_result172[24]^and_result172[25]^and_result172[26]^and_result172[27]^and_result172[28]^and_result172[29]^and_result172[30]^and_result172[31]^and_result172[32]^and_result172[33]^and_result172[34]^and_result172[35]^and_result172[36]^and_result172[37]^and_result172[38]^and_result172[39]^and_result172[40]^and_result172[41]^and_result172[42]^and_result172[43]^and_result172[44]^and_result172[45]^and_result172[46]^and_result172[47]^and_result172[48]^and_result172[49]^and_result172[50]^and_result172[51]^and_result172[52]^and_result172[53]^and_result172[54]^and_result172[55]^and_result172[56]^and_result172[57]^and_result172[58]^and_result172[59]^and_result172[60]^and_result172[61]^and_result172[62]^and_result172[63]^and_result172[64]^and_result172[65]^and_result172[66]^and_result172[67]^and_result172[68]^and_result172[69]^and_result172[70]^and_result172[71]^and_result172[72]^and_result172[73]^and_result172[74]^and_result172[75]^and_result172[76]^and_result172[77]^and_result172[78]^and_result172[79]^and_result172[80]^and_result172[81]^and_result172[82]^and_result172[83]^and_result172[84]^and_result172[85]^and_result172[86]^and_result172[87]^and_result172[88]^and_result172[89]^and_result172[90]^and_result172[91]^and_result172[92]^and_result172[93]^and_result172[94]^and_result172[95]^and_result172[96]^and_result172[97]^and_result172[98]^and_result172[99]^and_result172[100]^and_result172[101]^and_result172[102]^and_result172[103]^and_result172[104]^and_result172[105]^and_result172[106]^and_result172[107]^and_result172[108]^and_result172[109]^and_result172[110]^and_result172[111]^and_result172[112]^and_result172[113]^and_result172[114]^and_result172[115]^and_result172[116]^and_result172[117]^and_result172[118]^and_result172[119]^and_result172[120]^and_result172[121]^and_result172[122]^and_result172[123]^and_result172[124]^and_result172[125]^and_result172[126]^and_result172[127]^and_result172[128]^and_result172[129]^and_result172[130]^and_result172[131]^and_result172[132]^and_result172[133]^and_result172[134]^and_result172[135]^and_result172[136]^and_result172[137]^and_result172[138]^and_result172[139]^and_result172[140]^and_result172[141]^and_result172[142]^and_result172[143]^and_result172[144]^and_result172[145]^and_result172[146]^and_result172[147]^and_result172[148]^and_result172[149]^and_result172[150]^and_result172[151]^and_result172[152]^and_result172[153]^and_result172[154]^and_result172[155]^and_result172[156]^and_result172[157]^and_result172[158]^and_result172[159]^and_result172[160]^and_result172[161]^and_result172[162]^and_result172[163]^and_result172[164]^and_result172[165]^and_result172[166]^and_result172[167]^and_result172[168]^and_result172[169]^and_result172[170]^and_result172[171]^and_result172[172]^and_result172[173]^and_result172[174]^and_result172[175]^and_result172[176]^and_result172[177]^and_result172[178]^and_result172[179]^and_result172[180]^and_result172[181]^and_result172[182]^and_result172[183]^and_result172[184]^and_result172[185]^and_result172[186]^and_result172[187]^and_result172[188]^and_result172[189]^and_result172[190]^and_result172[191]^and_result172[192]^and_result172[193]^and_result172[194]^and_result172[195]^and_result172[196]^and_result172[197]^and_result172[198]^and_result172[199]^and_result172[200]^and_result172[201]^and_result172[202]^and_result172[203]^and_result172[204]^and_result172[205]^and_result172[206]^and_result172[207]^and_result172[208]^and_result172[209]^and_result172[210]^and_result172[211]^and_result172[212]^and_result172[213]^and_result172[214]^and_result172[215]^and_result172[216]^and_result172[217]^and_result172[218]^and_result172[219]^and_result172[220]^and_result172[221]^and_result172[222]^and_result172[223]^and_result172[224]^and_result172[225]^and_result172[226]^and_result172[227]^and_result172[228]^and_result172[229]^and_result172[230]^and_result172[231]^and_result172[232]^and_result172[233]^and_result172[234]^and_result172[235]^and_result172[236]^and_result172[237]^and_result172[238]^and_result172[239]^and_result172[240]^and_result172[241]^and_result172[242]^and_result172[243]^and_result172[244]^and_result172[245]^and_result172[246]^and_result172[247]^and_result172[248]^and_result172[249]^and_result172[250]^and_result172[251]^and_result172[252]^and_result172[253]^and_result172[254];
assign key[173]=and_result173[0]^and_result173[1]^and_result173[2]^and_result173[3]^and_result173[4]^and_result173[5]^and_result173[6]^and_result173[7]^and_result173[8]^and_result173[9]^and_result173[10]^and_result173[11]^and_result173[12]^and_result173[13]^and_result173[14]^and_result173[15]^and_result173[16]^and_result173[17]^and_result173[18]^and_result173[19]^and_result173[20]^and_result173[21]^and_result173[22]^and_result173[23]^and_result173[24]^and_result173[25]^and_result173[26]^and_result173[27]^and_result173[28]^and_result173[29]^and_result173[30]^and_result173[31]^and_result173[32]^and_result173[33]^and_result173[34]^and_result173[35]^and_result173[36]^and_result173[37]^and_result173[38]^and_result173[39]^and_result173[40]^and_result173[41]^and_result173[42]^and_result173[43]^and_result173[44]^and_result173[45]^and_result173[46]^and_result173[47]^and_result173[48]^and_result173[49]^and_result173[50]^and_result173[51]^and_result173[52]^and_result173[53]^and_result173[54]^and_result173[55]^and_result173[56]^and_result173[57]^and_result173[58]^and_result173[59]^and_result173[60]^and_result173[61]^and_result173[62]^and_result173[63]^and_result173[64]^and_result173[65]^and_result173[66]^and_result173[67]^and_result173[68]^and_result173[69]^and_result173[70]^and_result173[71]^and_result173[72]^and_result173[73]^and_result173[74]^and_result173[75]^and_result173[76]^and_result173[77]^and_result173[78]^and_result173[79]^and_result173[80]^and_result173[81]^and_result173[82]^and_result173[83]^and_result173[84]^and_result173[85]^and_result173[86]^and_result173[87]^and_result173[88]^and_result173[89]^and_result173[90]^and_result173[91]^and_result173[92]^and_result173[93]^and_result173[94]^and_result173[95]^and_result173[96]^and_result173[97]^and_result173[98]^and_result173[99]^and_result173[100]^and_result173[101]^and_result173[102]^and_result173[103]^and_result173[104]^and_result173[105]^and_result173[106]^and_result173[107]^and_result173[108]^and_result173[109]^and_result173[110]^and_result173[111]^and_result173[112]^and_result173[113]^and_result173[114]^and_result173[115]^and_result173[116]^and_result173[117]^and_result173[118]^and_result173[119]^and_result173[120]^and_result173[121]^and_result173[122]^and_result173[123]^and_result173[124]^and_result173[125]^and_result173[126]^and_result173[127]^and_result173[128]^and_result173[129]^and_result173[130]^and_result173[131]^and_result173[132]^and_result173[133]^and_result173[134]^and_result173[135]^and_result173[136]^and_result173[137]^and_result173[138]^and_result173[139]^and_result173[140]^and_result173[141]^and_result173[142]^and_result173[143]^and_result173[144]^and_result173[145]^and_result173[146]^and_result173[147]^and_result173[148]^and_result173[149]^and_result173[150]^and_result173[151]^and_result173[152]^and_result173[153]^and_result173[154]^and_result173[155]^and_result173[156]^and_result173[157]^and_result173[158]^and_result173[159]^and_result173[160]^and_result173[161]^and_result173[162]^and_result173[163]^and_result173[164]^and_result173[165]^and_result173[166]^and_result173[167]^and_result173[168]^and_result173[169]^and_result173[170]^and_result173[171]^and_result173[172]^and_result173[173]^and_result173[174]^and_result173[175]^and_result173[176]^and_result173[177]^and_result173[178]^and_result173[179]^and_result173[180]^and_result173[181]^and_result173[182]^and_result173[183]^and_result173[184]^and_result173[185]^and_result173[186]^and_result173[187]^and_result173[188]^and_result173[189]^and_result173[190]^and_result173[191]^and_result173[192]^and_result173[193]^and_result173[194]^and_result173[195]^and_result173[196]^and_result173[197]^and_result173[198]^and_result173[199]^and_result173[200]^and_result173[201]^and_result173[202]^and_result173[203]^and_result173[204]^and_result173[205]^and_result173[206]^and_result173[207]^and_result173[208]^and_result173[209]^and_result173[210]^and_result173[211]^and_result173[212]^and_result173[213]^and_result173[214]^and_result173[215]^and_result173[216]^and_result173[217]^and_result173[218]^and_result173[219]^and_result173[220]^and_result173[221]^and_result173[222]^and_result173[223]^and_result173[224]^and_result173[225]^and_result173[226]^and_result173[227]^and_result173[228]^and_result173[229]^and_result173[230]^and_result173[231]^and_result173[232]^and_result173[233]^and_result173[234]^and_result173[235]^and_result173[236]^and_result173[237]^and_result173[238]^and_result173[239]^and_result173[240]^and_result173[241]^and_result173[242]^and_result173[243]^and_result173[244]^and_result173[245]^and_result173[246]^and_result173[247]^and_result173[248]^and_result173[249]^and_result173[250]^and_result173[251]^and_result173[252]^and_result173[253]^and_result173[254];
assign key[174]=and_result174[0]^and_result174[1]^and_result174[2]^and_result174[3]^and_result174[4]^and_result174[5]^and_result174[6]^and_result174[7]^and_result174[8]^and_result174[9]^and_result174[10]^and_result174[11]^and_result174[12]^and_result174[13]^and_result174[14]^and_result174[15]^and_result174[16]^and_result174[17]^and_result174[18]^and_result174[19]^and_result174[20]^and_result174[21]^and_result174[22]^and_result174[23]^and_result174[24]^and_result174[25]^and_result174[26]^and_result174[27]^and_result174[28]^and_result174[29]^and_result174[30]^and_result174[31]^and_result174[32]^and_result174[33]^and_result174[34]^and_result174[35]^and_result174[36]^and_result174[37]^and_result174[38]^and_result174[39]^and_result174[40]^and_result174[41]^and_result174[42]^and_result174[43]^and_result174[44]^and_result174[45]^and_result174[46]^and_result174[47]^and_result174[48]^and_result174[49]^and_result174[50]^and_result174[51]^and_result174[52]^and_result174[53]^and_result174[54]^and_result174[55]^and_result174[56]^and_result174[57]^and_result174[58]^and_result174[59]^and_result174[60]^and_result174[61]^and_result174[62]^and_result174[63]^and_result174[64]^and_result174[65]^and_result174[66]^and_result174[67]^and_result174[68]^and_result174[69]^and_result174[70]^and_result174[71]^and_result174[72]^and_result174[73]^and_result174[74]^and_result174[75]^and_result174[76]^and_result174[77]^and_result174[78]^and_result174[79]^and_result174[80]^and_result174[81]^and_result174[82]^and_result174[83]^and_result174[84]^and_result174[85]^and_result174[86]^and_result174[87]^and_result174[88]^and_result174[89]^and_result174[90]^and_result174[91]^and_result174[92]^and_result174[93]^and_result174[94]^and_result174[95]^and_result174[96]^and_result174[97]^and_result174[98]^and_result174[99]^and_result174[100]^and_result174[101]^and_result174[102]^and_result174[103]^and_result174[104]^and_result174[105]^and_result174[106]^and_result174[107]^and_result174[108]^and_result174[109]^and_result174[110]^and_result174[111]^and_result174[112]^and_result174[113]^and_result174[114]^and_result174[115]^and_result174[116]^and_result174[117]^and_result174[118]^and_result174[119]^and_result174[120]^and_result174[121]^and_result174[122]^and_result174[123]^and_result174[124]^and_result174[125]^and_result174[126]^and_result174[127]^and_result174[128]^and_result174[129]^and_result174[130]^and_result174[131]^and_result174[132]^and_result174[133]^and_result174[134]^and_result174[135]^and_result174[136]^and_result174[137]^and_result174[138]^and_result174[139]^and_result174[140]^and_result174[141]^and_result174[142]^and_result174[143]^and_result174[144]^and_result174[145]^and_result174[146]^and_result174[147]^and_result174[148]^and_result174[149]^and_result174[150]^and_result174[151]^and_result174[152]^and_result174[153]^and_result174[154]^and_result174[155]^and_result174[156]^and_result174[157]^and_result174[158]^and_result174[159]^and_result174[160]^and_result174[161]^and_result174[162]^and_result174[163]^and_result174[164]^and_result174[165]^and_result174[166]^and_result174[167]^and_result174[168]^and_result174[169]^and_result174[170]^and_result174[171]^and_result174[172]^and_result174[173]^and_result174[174]^and_result174[175]^and_result174[176]^and_result174[177]^and_result174[178]^and_result174[179]^and_result174[180]^and_result174[181]^and_result174[182]^and_result174[183]^and_result174[184]^and_result174[185]^and_result174[186]^and_result174[187]^and_result174[188]^and_result174[189]^and_result174[190]^and_result174[191]^and_result174[192]^and_result174[193]^and_result174[194]^and_result174[195]^and_result174[196]^and_result174[197]^and_result174[198]^and_result174[199]^and_result174[200]^and_result174[201]^and_result174[202]^and_result174[203]^and_result174[204]^and_result174[205]^and_result174[206]^and_result174[207]^and_result174[208]^and_result174[209]^and_result174[210]^and_result174[211]^and_result174[212]^and_result174[213]^and_result174[214]^and_result174[215]^and_result174[216]^and_result174[217]^and_result174[218]^and_result174[219]^and_result174[220]^and_result174[221]^and_result174[222]^and_result174[223]^and_result174[224]^and_result174[225]^and_result174[226]^and_result174[227]^and_result174[228]^and_result174[229]^and_result174[230]^and_result174[231]^and_result174[232]^and_result174[233]^and_result174[234]^and_result174[235]^and_result174[236]^and_result174[237]^and_result174[238]^and_result174[239]^and_result174[240]^and_result174[241]^and_result174[242]^and_result174[243]^and_result174[244]^and_result174[245]^and_result174[246]^and_result174[247]^and_result174[248]^and_result174[249]^and_result174[250]^and_result174[251]^and_result174[252]^and_result174[253]^and_result174[254];
assign key[175]=and_result175[0]^and_result175[1]^and_result175[2]^and_result175[3]^and_result175[4]^and_result175[5]^and_result175[6]^and_result175[7]^and_result175[8]^and_result175[9]^and_result175[10]^and_result175[11]^and_result175[12]^and_result175[13]^and_result175[14]^and_result175[15]^and_result175[16]^and_result175[17]^and_result175[18]^and_result175[19]^and_result175[20]^and_result175[21]^and_result175[22]^and_result175[23]^and_result175[24]^and_result175[25]^and_result175[26]^and_result175[27]^and_result175[28]^and_result175[29]^and_result175[30]^and_result175[31]^and_result175[32]^and_result175[33]^and_result175[34]^and_result175[35]^and_result175[36]^and_result175[37]^and_result175[38]^and_result175[39]^and_result175[40]^and_result175[41]^and_result175[42]^and_result175[43]^and_result175[44]^and_result175[45]^and_result175[46]^and_result175[47]^and_result175[48]^and_result175[49]^and_result175[50]^and_result175[51]^and_result175[52]^and_result175[53]^and_result175[54]^and_result175[55]^and_result175[56]^and_result175[57]^and_result175[58]^and_result175[59]^and_result175[60]^and_result175[61]^and_result175[62]^and_result175[63]^and_result175[64]^and_result175[65]^and_result175[66]^and_result175[67]^and_result175[68]^and_result175[69]^and_result175[70]^and_result175[71]^and_result175[72]^and_result175[73]^and_result175[74]^and_result175[75]^and_result175[76]^and_result175[77]^and_result175[78]^and_result175[79]^and_result175[80]^and_result175[81]^and_result175[82]^and_result175[83]^and_result175[84]^and_result175[85]^and_result175[86]^and_result175[87]^and_result175[88]^and_result175[89]^and_result175[90]^and_result175[91]^and_result175[92]^and_result175[93]^and_result175[94]^and_result175[95]^and_result175[96]^and_result175[97]^and_result175[98]^and_result175[99]^and_result175[100]^and_result175[101]^and_result175[102]^and_result175[103]^and_result175[104]^and_result175[105]^and_result175[106]^and_result175[107]^and_result175[108]^and_result175[109]^and_result175[110]^and_result175[111]^and_result175[112]^and_result175[113]^and_result175[114]^and_result175[115]^and_result175[116]^and_result175[117]^and_result175[118]^and_result175[119]^and_result175[120]^and_result175[121]^and_result175[122]^and_result175[123]^and_result175[124]^and_result175[125]^and_result175[126]^and_result175[127]^and_result175[128]^and_result175[129]^and_result175[130]^and_result175[131]^and_result175[132]^and_result175[133]^and_result175[134]^and_result175[135]^and_result175[136]^and_result175[137]^and_result175[138]^and_result175[139]^and_result175[140]^and_result175[141]^and_result175[142]^and_result175[143]^and_result175[144]^and_result175[145]^and_result175[146]^and_result175[147]^and_result175[148]^and_result175[149]^and_result175[150]^and_result175[151]^and_result175[152]^and_result175[153]^and_result175[154]^and_result175[155]^and_result175[156]^and_result175[157]^and_result175[158]^and_result175[159]^and_result175[160]^and_result175[161]^and_result175[162]^and_result175[163]^and_result175[164]^and_result175[165]^and_result175[166]^and_result175[167]^and_result175[168]^and_result175[169]^and_result175[170]^and_result175[171]^and_result175[172]^and_result175[173]^and_result175[174]^and_result175[175]^and_result175[176]^and_result175[177]^and_result175[178]^and_result175[179]^and_result175[180]^and_result175[181]^and_result175[182]^and_result175[183]^and_result175[184]^and_result175[185]^and_result175[186]^and_result175[187]^and_result175[188]^and_result175[189]^and_result175[190]^and_result175[191]^and_result175[192]^and_result175[193]^and_result175[194]^and_result175[195]^and_result175[196]^and_result175[197]^and_result175[198]^and_result175[199]^and_result175[200]^and_result175[201]^and_result175[202]^and_result175[203]^and_result175[204]^and_result175[205]^and_result175[206]^and_result175[207]^and_result175[208]^and_result175[209]^and_result175[210]^and_result175[211]^and_result175[212]^and_result175[213]^and_result175[214]^and_result175[215]^and_result175[216]^and_result175[217]^and_result175[218]^and_result175[219]^and_result175[220]^and_result175[221]^and_result175[222]^and_result175[223]^and_result175[224]^and_result175[225]^and_result175[226]^and_result175[227]^and_result175[228]^and_result175[229]^and_result175[230]^and_result175[231]^and_result175[232]^and_result175[233]^and_result175[234]^and_result175[235]^and_result175[236]^and_result175[237]^and_result175[238]^and_result175[239]^and_result175[240]^and_result175[241]^and_result175[242]^and_result175[243]^and_result175[244]^and_result175[245]^and_result175[246]^and_result175[247]^and_result175[248]^and_result175[249]^and_result175[250]^and_result175[251]^and_result175[252]^and_result175[253]^and_result175[254];
assign key[176]=and_result176[0]^and_result176[1]^and_result176[2]^and_result176[3]^and_result176[4]^and_result176[5]^and_result176[6]^and_result176[7]^and_result176[8]^and_result176[9]^and_result176[10]^and_result176[11]^and_result176[12]^and_result176[13]^and_result176[14]^and_result176[15]^and_result176[16]^and_result176[17]^and_result176[18]^and_result176[19]^and_result176[20]^and_result176[21]^and_result176[22]^and_result176[23]^and_result176[24]^and_result176[25]^and_result176[26]^and_result176[27]^and_result176[28]^and_result176[29]^and_result176[30]^and_result176[31]^and_result176[32]^and_result176[33]^and_result176[34]^and_result176[35]^and_result176[36]^and_result176[37]^and_result176[38]^and_result176[39]^and_result176[40]^and_result176[41]^and_result176[42]^and_result176[43]^and_result176[44]^and_result176[45]^and_result176[46]^and_result176[47]^and_result176[48]^and_result176[49]^and_result176[50]^and_result176[51]^and_result176[52]^and_result176[53]^and_result176[54]^and_result176[55]^and_result176[56]^and_result176[57]^and_result176[58]^and_result176[59]^and_result176[60]^and_result176[61]^and_result176[62]^and_result176[63]^and_result176[64]^and_result176[65]^and_result176[66]^and_result176[67]^and_result176[68]^and_result176[69]^and_result176[70]^and_result176[71]^and_result176[72]^and_result176[73]^and_result176[74]^and_result176[75]^and_result176[76]^and_result176[77]^and_result176[78]^and_result176[79]^and_result176[80]^and_result176[81]^and_result176[82]^and_result176[83]^and_result176[84]^and_result176[85]^and_result176[86]^and_result176[87]^and_result176[88]^and_result176[89]^and_result176[90]^and_result176[91]^and_result176[92]^and_result176[93]^and_result176[94]^and_result176[95]^and_result176[96]^and_result176[97]^and_result176[98]^and_result176[99]^and_result176[100]^and_result176[101]^and_result176[102]^and_result176[103]^and_result176[104]^and_result176[105]^and_result176[106]^and_result176[107]^and_result176[108]^and_result176[109]^and_result176[110]^and_result176[111]^and_result176[112]^and_result176[113]^and_result176[114]^and_result176[115]^and_result176[116]^and_result176[117]^and_result176[118]^and_result176[119]^and_result176[120]^and_result176[121]^and_result176[122]^and_result176[123]^and_result176[124]^and_result176[125]^and_result176[126]^and_result176[127]^and_result176[128]^and_result176[129]^and_result176[130]^and_result176[131]^and_result176[132]^and_result176[133]^and_result176[134]^and_result176[135]^and_result176[136]^and_result176[137]^and_result176[138]^and_result176[139]^and_result176[140]^and_result176[141]^and_result176[142]^and_result176[143]^and_result176[144]^and_result176[145]^and_result176[146]^and_result176[147]^and_result176[148]^and_result176[149]^and_result176[150]^and_result176[151]^and_result176[152]^and_result176[153]^and_result176[154]^and_result176[155]^and_result176[156]^and_result176[157]^and_result176[158]^and_result176[159]^and_result176[160]^and_result176[161]^and_result176[162]^and_result176[163]^and_result176[164]^and_result176[165]^and_result176[166]^and_result176[167]^and_result176[168]^and_result176[169]^and_result176[170]^and_result176[171]^and_result176[172]^and_result176[173]^and_result176[174]^and_result176[175]^and_result176[176]^and_result176[177]^and_result176[178]^and_result176[179]^and_result176[180]^and_result176[181]^and_result176[182]^and_result176[183]^and_result176[184]^and_result176[185]^and_result176[186]^and_result176[187]^and_result176[188]^and_result176[189]^and_result176[190]^and_result176[191]^and_result176[192]^and_result176[193]^and_result176[194]^and_result176[195]^and_result176[196]^and_result176[197]^and_result176[198]^and_result176[199]^and_result176[200]^and_result176[201]^and_result176[202]^and_result176[203]^and_result176[204]^and_result176[205]^and_result176[206]^and_result176[207]^and_result176[208]^and_result176[209]^and_result176[210]^and_result176[211]^and_result176[212]^and_result176[213]^and_result176[214]^and_result176[215]^and_result176[216]^and_result176[217]^and_result176[218]^and_result176[219]^and_result176[220]^and_result176[221]^and_result176[222]^and_result176[223]^and_result176[224]^and_result176[225]^and_result176[226]^and_result176[227]^and_result176[228]^and_result176[229]^and_result176[230]^and_result176[231]^and_result176[232]^and_result176[233]^and_result176[234]^and_result176[235]^and_result176[236]^and_result176[237]^and_result176[238]^and_result176[239]^and_result176[240]^and_result176[241]^and_result176[242]^and_result176[243]^and_result176[244]^and_result176[245]^and_result176[246]^and_result176[247]^and_result176[248]^and_result176[249]^and_result176[250]^and_result176[251]^and_result176[252]^and_result176[253]^and_result176[254];
assign key[177]=and_result177[0]^and_result177[1]^and_result177[2]^and_result177[3]^and_result177[4]^and_result177[5]^and_result177[6]^and_result177[7]^and_result177[8]^and_result177[9]^and_result177[10]^and_result177[11]^and_result177[12]^and_result177[13]^and_result177[14]^and_result177[15]^and_result177[16]^and_result177[17]^and_result177[18]^and_result177[19]^and_result177[20]^and_result177[21]^and_result177[22]^and_result177[23]^and_result177[24]^and_result177[25]^and_result177[26]^and_result177[27]^and_result177[28]^and_result177[29]^and_result177[30]^and_result177[31]^and_result177[32]^and_result177[33]^and_result177[34]^and_result177[35]^and_result177[36]^and_result177[37]^and_result177[38]^and_result177[39]^and_result177[40]^and_result177[41]^and_result177[42]^and_result177[43]^and_result177[44]^and_result177[45]^and_result177[46]^and_result177[47]^and_result177[48]^and_result177[49]^and_result177[50]^and_result177[51]^and_result177[52]^and_result177[53]^and_result177[54]^and_result177[55]^and_result177[56]^and_result177[57]^and_result177[58]^and_result177[59]^and_result177[60]^and_result177[61]^and_result177[62]^and_result177[63]^and_result177[64]^and_result177[65]^and_result177[66]^and_result177[67]^and_result177[68]^and_result177[69]^and_result177[70]^and_result177[71]^and_result177[72]^and_result177[73]^and_result177[74]^and_result177[75]^and_result177[76]^and_result177[77]^and_result177[78]^and_result177[79]^and_result177[80]^and_result177[81]^and_result177[82]^and_result177[83]^and_result177[84]^and_result177[85]^and_result177[86]^and_result177[87]^and_result177[88]^and_result177[89]^and_result177[90]^and_result177[91]^and_result177[92]^and_result177[93]^and_result177[94]^and_result177[95]^and_result177[96]^and_result177[97]^and_result177[98]^and_result177[99]^and_result177[100]^and_result177[101]^and_result177[102]^and_result177[103]^and_result177[104]^and_result177[105]^and_result177[106]^and_result177[107]^and_result177[108]^and_result177[109]^and_result177[110]^and_result177[111]^and_result177[112]^and_result177[113]^and_result177[114]^and_result177[115]^and_result177[116]^and_result177[117]^and_result177[118]^and_result177[119]^and_result177[120]^and_result177[121]^and_result177[122]^and_result177[123]^and_result177[124]^and_result177[125]^and_result177[126]^and_result177[127]^and_result177[128]^and_result177[129]^and_result177[130]^and_result177[131]^and_result177[132]^and_result177[133]^and_result177[134]^and_result177[135]^and_result177[136]^and_result177[137]^and_result177[138]^and_result177[139]^and_result177[140]^and_result177[141]^and_result177[142]^and_result177[143]^and_result177[144]^and_result177[145]^and_result177[146]^and_result177[147]^and_result177[148]^and_result177[149]^and_result177[150]^and_result177[151]^and_result177[152]^and_result177[153]^and_result177[154]^and_result177[155]^and_result177[156]^and_result177[157]^and_result177[158]^and_result177[159]^and_result177[160]^and_result177[161]^and_result177[162]^and_result177[163]^and_result177[164]^and_result177[165]^and_result177[166]^and_result177[167]^and_result177[168]^and_result177[169]^and_result177[170]^and_result177[171]^and_result177[172]^and_result177[173]^and_result177[174]^and_result177[175]^and_result177[176]^and_result177[177]^and_result177[178]^and_result177[179]^and_result177[180]^and_result177[181]^and_result177[182]^and_result177[183]^and_result177[184]^and_result177[185]^and_result177[186]^and_result177[187]^and_result177[188]^and_result177[189]^and_result177[190]^and_result177[191]^and_result177[192]^and_result177[193]^and_result177[194]^and_result177[195]^and_result177[196]^and_result177[197]^and_result177[198]^and_result177[199]^and_result177[200]^and_result177[201]^and_result177[202]^and_result177[203]^and_result177[204]^and_result177[205]^and_result177[206]^and_result177[207]^and_result177[208]^and_result177[209]^and_result177[210]^and_result177[211]^and_result177[212]^and_result177[213]^and_result177[214]^and_result177[215]^and_result177[216]^and_result177[217]^and_result177[218]^and_result177[219]^and_result177[220]^and_result177[221]^and_result177[222]^and_result177[223]^and_result177[224]^and_result177[225]^and_result177[226]^and_result177[227]^and_result177[228]^and_result177[229]^and_result177[230]^and_result177[231]^and_result177[232]^and_result177[233]^and_result177[234]^and_result177[235]^and_result177[236]^and_result177[237]^and_result177[238]^and_result177[239]^and_result177[240]^and_result177[241]^and_result177[242]^and_result177[243]^and_result177[244]^and_result177[245]^and_result177[246]^and_result177[247]^and_result177[248]^and_result177[249]^and_result177[250]^and_result177[251]^and_result177[252]^and_result177[253]^and_result177[254];
assign key[178]=and_result178[0]^and_result178[1]^and_result178[2]^and_result178[3]^and_result178[4]^and_result178[5]^and_result178[6]^and_result178[7]^and_result178[8]^and_result178[9]^and_result178[10]^and_result178[11]^and_result178[12]^and_result178[13]^and_result178[14]^and_result178[15]^and_result178[16]^and_result178[17]^and_result178[18]^and_result178[19]^and_result178[20]^and_result178[21]^and_result178[22]^and_result178[23]^and_result178[24]^and_result178[25]^and_result178[26]^and_result178[27]^and_result178[28]^and_result178[29]^and_result178[30]^and_result178[31]^and_result178[32]^and_result178[33]^and_result178[34]^and_result178[35]^and_result178[36]^and_result178[37]^and_result178[38]^and_result178[39]^and_result178[40]^and_result178[41]^and_result178[42]^and_result178[43]^and_result178[44]^and_result178[45]^and_result178[46]^and_result178[47]^and_result178[48]^and_result178[49]^and_result178[50]^and_result178[51]^and_result178[52]^and_result178[53]^and_result178[54]^and_result178[55]^and_result178[56]^and_result178[57]^and_result178[58]^and_result178[59]^and_result178[60]^and_result178[61]^and_result178[62]^and_result178[63]^and_result178[64]^and_result178[65]^and_result178[66]^and_result178[67]^and_result178[68]^and_result178[69]^and_result178[70]^and_result178[71]^and_result178[72]^and_result178[73]^and_result178[74]^and_result178[75]^and_result178[76]^and_result178[77]^and_result178[78]^and_result178[79]^and_result178[80]^and_result178[81]^and_result178[82]^and_result178[83]^and_result178[84]^and_result178[85]^and_result178[86]^and_result178[87]^and_result178[88]^and_result178[89]^and_result178[90]^and_result178[91]^and_result178[92]^and_result178[93]^and_result178[94]^and_result178[95]^and_result178[96]^and_result178[97]^and_result178[98]^and_result178[99]^and_result178[100]^and_result178[101]^and_result178[102]^and_result178[103]^and_result178[104]^and_result178[105]^and_result178[106]^and_result178[107]^and_result178[108]^and_result178[109]^and_result178[110]^and_result178[111]^and_result178[112]^and_result178[113]^and_result178[114]^and_result178[115]^and_result178[116]^and_result178[117]^and_result178[118]^and_result178[119]^and_result178[120]^and_result178[121]^and_result178[122]^and_result178[123]^and_result178[124]^and_result178[125]^and_result178[126]^and_result178[127]^and_result178[128]^and_result178[129]^and_result178[130]^and_result178[131]^and_result178[132]^and_result178[133]^and_result178[134]^and_result178[135]^and_result178[136]^and_result178[137]^and_result178[138]^and_result178[139]^and_result178[140]^and_result178[141]^and_result178[142]^and_result178[143]^and_result178[144]^and_result178[145]^and_result178[146]^and_result178[147]^and_result178[148]^and_result178[149]^and_result178[150]^and_result178[151]^and_result178[152]^and_result178[153]^and_result178[154]^and_result178[155]^and_result178[156]^and_result178[157]^and_result178[158]^and_result178[159]^and_result178[160]^and_result178[161]^and_result178[162]^and_result178[163]^and_result178[164]^and_result178[165]^and_result178[166]^and_result178[167]^and_result178[168]^and_result178[169]^and_result178[170]^and_result178[171]^and_result178[172]^and_result178[173]^and_result178[174]^and_result178[175]^and_result178[176]^and_result178[177]^and_result178[178]^and_result178[179]^and_result178[180]^and_result178[181]^and_result178[182]^and_result178[183]^and_result178[184]^and_result178[185]^and_result178[186]^and_result178[187]^and_result178[188]^and_result178[189]^and_result178[190]^and_result178[191]^and_result178[192]^and_result178[193]^and_result178[194]^and_result178[195]^and_result178[196]^and_result178[197]^and_result178[198]^and_result178[199]^and_result178[200]^and_result178[201]^and_result178[202]^and_result178[203]^and_result178[204]^and_result178[205]^and_result178[206]^and_result178[207]^and_result178[208]^and_result178[209]^and_result178[210]^and_result178[211]^and_result178[212]^and_result178[213]^and_result178[214]^and_result178[215]^and_result178[216]^and_result178[217]^and_result178[218]^and_result178[219]^and_result178[220]^and_result178[221]^and_result178[222]^and_result178[223]^and_result178[224]^and_result178[225]^and_result178[226]^and_result178[227]^and_result178[228]^and_result178[229]^and_result178[230]^and_result178[231]^and_result178[232]^and_result178[233]^and_result178[234]^and_result178[235]^and_result178[236]^and_result178[237]^and_result178[238]^and_result178[239]^and_result178[240]^and_result178[241]^and_result178[242]^and_result178[243]^and_result178[244]^and_result178[245]^and_result178[246]^and_result178[247]^and_result178[248]^and_result178[249]^and_result178[250]^and_result178[251]^and_result178[252]^and_result178[253]^and_result178[254];
assign key[179]=and_result179[0]^and_result179[1]^and_result179[2]^and_result179[3]^and_result179[4]^and_result179[5]^and_result179[6]^and_result179[7]^and_result179[8]^and_result179[9]^and_result179[10]^and_result179[11]^and_result179[12]^and_result179[13]^and_result179[14]^and_result179[15]^and_result179[16]^and_result179[17]^and_result179[18]^and_result179[19]^and_result179[20]^and_result179[21]^and_result179[22]^and_result179[23]^and_result179[24]^and_result179[25]^and_result179[26]^and_result179[27]^and_result179[28]^and_result179[29]^and_result179[30]^and_result179[31]^and_result179[32]^and_result179[33]^and_result179[34]^and_result179[35]^and_result179[36]^and_result179[37]^and_result179[38]^and_result179[39]^and_result179[40]^and_result179[41]^and_result179[42]^and_result179[43]^and_result179[44]^and_result179[45]^and_result179[46]^and_result179[47]^and_result179[48]^and_result179[49]^and_result179[50]^and_result179[51]^and_result179[52]^and_result179[53]^and_result179[54]^and_result179[55]^and_result179[56]^and_result179[57]^and_result179[58]^and_result179[59]^and_result179[60]^and_result179[61]^and_result179[62]^and_result179[63]^and_result179[64]^and_result179[65]^and_result179[66]^and_result179[67]^and_result179[68]^and_result179[69]^and_result179[70]^and_result179[71]^and_result179[72]^and_result179[73]^and_result179[74]^and_result179[75]^and_result179[76]^and_result179[77]^and_result179[78]^and_result179[79]^and_result179[80]^and_result179[81]^and_result179[82]^and_result179[83]^and_result179[84]^and_result179[85]^and_result179[86]^and_result179[87]^and_result179[88]^and_result179[89]^and_result179[90]^and_result179[91]^and_result179[92]^and_result179[93]^and_result179[94]^and_result179[95]^and_result179[96]^and_result179[97]^and_result179[98]^and_result179[99]^and_result179[100]^and_result179[101]^and_result179[102]^and_result179[103]^and_result179[104]^and_result179[105]^and_result179[106]^and_result179[107]^and_result179[108]^and_result179[109]^and_result179[110]^and_result179[111]^and_result179[112]^and_result179[113]^and_result179[114]^and_result179[115]^and_result179[116]^and_result179[117]^and_result179[118]^and_result179[119]^and_result179[120]^and_result179[121]^and_result179[122]^and_result179[123]^and_result179[124]^and_result179[125]^and_result179[126]^and_result179[127]^and_result179[128]^and_result179[129]^and_result179[130]^and_result179[131]^and_result179[132]^and_result179[133]^and_result179[134]^and_result179[135]^and_result179[136]^and_result179[137]^and_result179[138]^and_result179[139]^and_result179[140]^and_result179[141]^and_result179[142]^and_result179[143]^and_result179[144]^and_result179[145]^and_result179[146]^and_result179[147]^and_result179[148]^and_result179[149]^and_result179[150]^and_result179[151]^and_result179[152]^and_result179[153]^and_result179[154]^and_result179[155]^and_result179[156]^and_result179[157]^and_result179[158]^and_result179[159]^and_result179[160]^and_result179[161]^and_result179[162]^and_result179[163]^and_result179[164]^and_result179[165]^and_result179[166]^and_result179[167]^and_result179[168]^and_result179[169]^and_result179[170]^and_result179[171]^and_result179[172]^and_result179[173]^and_result179[174]^and_result179[175]^and_result179[176]^and_result179[177]^and_result179[178]^and_result179[179]^and_result179[180]^and_result179[181]^and_result179[182]^and_result179[183]^and_result179[184]^and_result179[185]^and_result179[186]^and_result179[187]^and_result179[188]^and_result179[189]^and_result179[190]^and_result179[191]^and_result179[192]^and_result179[193]^and_result179[194]^and_result179[195]^and_result179[196]^and_result179[197]^and_result179[198]^and_result179[199]^and_result179[200]^and_result179[201]^and_result179[202]^and_result179[203]^and_result179[204]^and_result179[205]^and_result179[206]^and_result179[207]^and_result179[208]^and_result179[209]^and_result179[210]^and_result179[211]^and_result179[212]^and_result179[213]^and_result179[214]^and_result179[215]^and_result179[216]^and_result179[217]^and_result179[218]^and_result179[219]^and_result179[220]^and_result179[221]^and_result179[222]^and_result179[223]^and_result179[224]^and_result179[225]^and_result179[226]^and_result179[227]^and_result179[228]^and_result179[229]^and_result179[230]^and_result179[231]^and_result179[232]^and_result179[233]^and_result179[234]^and_result179[235]^and_result179[236]^and_result179[237]^and_result179[238]^and_result179[239]^and_result179[240]^and_result179[241]^and_result179[242]^and_result179[243]^and_result179[244]^and_result179[245]^and_result179[246]^and_result179[247]^and_result179[248]^and_result179[249]^and_result179[250]^and_result179[251]^and_result179[252]^and_result179[253]^and_result179[254];
assign key[180]=and_result180[0]^and_result180[1]^and_result180[2]^and_result180[3]^and_result180[4]^and_result180[5]^and_result180[6]^and_result180[7]^and_result180[8]^and_result180[9]^and_result180[10]^and_result180[11]^and_result180[12]^and_result180[13]^and_result180[14]^and_result180[15]^and_result180[16]^and_result180[17]^and_result180[18]^and_result180[19]^and_result180[20]^and_result180[21]^and_result180[22]^and_result180[23]^and_result180[24]^and_result180[25]^and_result180[26]^and_result180[27]^and_result180[28]^and_result180[29]^and_result180[30]^and_result180[31]^and_result180[32]^and_result180[33]^and_result180[34]^and_result180[35]^and_result180[36]^and_result180[37]^and_result180[38]^and_result180[39]^and_result180[40]^and_result180[41]^and_result180[42]^and_result180[43]^and_result180[44]^and_result180[45]^and_result180[46]^and_result180[47]^and_result180[48]^and_result180[49]^and_result180[50]^and_result180[51]^and_result180[52]^and_result180[53]^and_result180[54]^and_result180[55]^and_result180[56]^and_result180[57]^and_result180[58]^and_result180[59]^and_result180[60]^and_result180[61]^and_result180[62]^and_result180[63]^and_result180[64]^and_result180[65]^and_result180[66]^and_result180[67]^and_result180[68]^and_result180[69]^and_result180[70]^and_result180[71]^and_result180[72]^and_result180[73]^and_result180[74]^and_result180[75]^and_result180[76]^and_result180[77]^and_result180[78]^and_result180[79]^and_result180[80]^and_result180[81]^and_result180[82]^and_result180[83]^and_result180[84]^and_result180[85]^and_result180[86]^and_result180[87]^and_result180[88]^and_result180[89]^and_result180[90]^and_result180[91]^and_result180[92]^and_result180[93]^and_result180[94]^and_result180[95]^and_result180[96]^and_result180[97]^and_result180[98]^and_result180[99]^and_result180[100]^and_result180[101]^and_result180[102]^and_result180[103]^and_result180[104]^and_result180[105]^and_result180[106]^and_result180[107]^and_result180[108]^and_result180[109]^and_result180[110]^and_result180[111]^and_result180[112]^and_result180[113]^and_result180[114]^and_result180[115]^and_result180[116]^and_result180[117]^and_result180[118]^and_result180[119]^and_result180[120]^and_result180[121]^and_result180[122]^and_result180[123]^and_result180[124]^and_result180[125]^and_result180[126]^and_result180[127]^and_result180[128]^and_result180[129]^and_result180[130]^and_result180[131]^and_result180[132]^and_result180[133]^and_result180[134]^and_result180[135]^and_result180[136]^and_result180[137]^and_result180[138]^and_result180[139]^and_result180[140]^and_result180[141]^and_result180[142]^and_result180[143]^and_result180[144]^and_result180[145]^and_result180[146]^and_result180[147]^and_result180[148]^and_result180[149]^and_result180[150]^and_result180[151]^and_result180[152]^and_result180[153]^and_result180[154]^and_result180[155]^and_result180[156]^and_result180[157]^and_result180[158]^and_result180[159]^and_result180[160]^and_result180[161]^and_result180[162]^and_result180[163]^and_result180[164]^and_result180[165]^and_result180[166]^and_result180[167]^and_result180[168]^and_result180[169]^and_result180[170]^and_result180[171]^and_result180[172]^and_result180[173]^and_result180[174]^and_result180[175]^and_result180[176]^and_result180[177]^and_result180[178]^and_result180[179]^and_result180[180]^and_result180[181]^and_result180[182]^and_result180[183]^and_result180[184]^and_result180[185]^and_result180[186]^and_result180[187]^and_result180[188]^and_result180[189]^and_result180[190]^and_result180[191]^and_result180[192]^and_result180[193]^and_result180[194]^and_result180[195]^and_result180[196]^and_result180[197]^and_result180[198]^and_result180[199]^and_result180[200]^and_result180[201]^and_result180[202]^and_result180[203]^and_result180[204]^and_result180[205]^and_result180[206]^and_result180[207]^and_result180[208]^and_result180[209]^and_result180[210]^and_result180[211]^and_result180[212]^and_result180[213]^and_result180[214]^and_result180[215]^and_result180[216]^and_result180[217]^and_result180[218]^and_result180[219]^and_result180[220]^and_result180[221]^and_result180[222]^and_result180[223]^and_result180[224]^and_result180[225]^and_result180[226]^and_result180[227]^and_result180[228]^and_result180[229]^and_result180[230]^and_result180[231]^and_result180[232]^and_result180[233]^and_result180[234]^and_result180[235]^and_result180[236]^and_result180[237]^and_result180[238]^and_result180[239]^and_result180[240]^and_result180[241]^and_result180[242]^and_result180[243]^and_result180[244]^and_result180[245]^and_result180[246]^and_result180[247]^and_result180[248]^and_result180[249]^and_result180[250]^and_result180[251]^and_result180[252]^and_result180[253]^and_result180[254];
assign key[181]=and_result181[0]^and_result181[1]^and_result181[2]^and_result181[3]^and_result181[4]^and_result181[5]^and_result181[6]^and_result181[7]^and_result181[8]^and_result181[9]^and_result181[10]^and_result181[11]^and_result181[12]^and_result181[13]^and_result181[14]^and_result181[15]^and_result181[16]^and_result181[17]^and_result181[18]^and_result181[19]^and_result181[20]^and_result181[21]^and_result181[22]^and_result181[23]^and_result181[24]^and_result181[25]^and_result181[26]^and_result181[27]^and_result181[28]^and_result181[29]^and_result181[30]^and_result181[31]^and_result181[32]^and_result181[33]^and_result181[34]^and_result181[35]^and_result181[36]^and_result181[37]^and_result181[38]^and_result181[39]^and_result181[40]^and_result181[41]^and_result181[42]^and_result181[43]^and_result181[44]^and_result181[45]^and_result181[46]^and_result181[47]^and_result181[48]^and_result181[49]^and_result181[50]^and_result181[51]^and_result181[52]^and_result181[53]^and_result181[54]^and_result181[55]^and_result181[56]^and_result181[57]^and_result181[58]^and_result181[59]^and_result181[60]^and_result181[61]^and_result181[62]^and_result181[63]^and_result181[64]^and_result181[65]^and_result181[66]^and_result181[67]^and_result181[68]^and_result181[69]^and_result181[70]^and_result181[71]^and_result181[72]^and_result181[73]^and_result181[74]^and_result181[75]^and_result181[76]^and_result181[77]^and_result181[78]^and_result181[79]^and_result181[80]^and_result181[81]^and_result181[82]^and_result181[83]^and_result181[84]^and_result181[85]^and_result181[86]^and_result181[87]^and_result181[88]^and_result181[89]^and_result181[90]^and_result181[91]^and_result181[92]^and_result181[93]^and_result181[94]^and_result181[95]^and_result181[96]^and_result181[97]^and_result181[98]^and_result181[99]^and_result181[100]^and_result181[101]^and_result181[102]^and_result181[103]^and_result181[104]^and_result181[105]^and_result181[106]^and_result181[107]^and_result181[108]^and_result181[109]^and_result181[110]^and_result181[111]^and_result181[112]^and_result181[113]^and_result181[114]^and_result181[115]^and_result181[116]^and_result181[117]^and_result181[118]^and_result181[119]^and_result181[120]^and_result181[121]^and_result181[122]^and_result181[123]^and_result181[124]^and_result181[125]^and_result181[126]^and_result181[127]^and_result181[128]^and_result181[129]^and_result181[130]^and_result181[131]^and_result181[132]^and_result181[133]^and_result181[134]^and_result181[135]^and_result181[136]^and_result181[137]^and_result181[138]^and_result181[139]^and_result181[140]^and_result181[141]^and_result181[142]^and_result181[143]^and_result181[144]^and_result181[145]^and_result181[146]^and_result181[147]^and_result181[148]^and_result181[149]^and_result181[150]^and_result181[151]^and_result181[152]^and_result181[153]^and_result181[154]^and_result181[155]^and_result181[156]^and_result181[157]^and_result181[158]^and_result181[159]^and_result181[160]^and_result181[161]^and_result181[162]^and_result181[163]^and_result181[164]^and_result181[165]^and_result181[166]^and_result181[167]^and_result181[168]^and_result181[169]^and_result181[170]^and_result181[171]^and_result181[172]^and_result181[173]^and_result181[174]^and_result181[175]^and_result181[176]^and_result181[177]^and_result181[178]^and_result181[179]^and_result181[180]^and_result181[181]^and_result181[182]^and_result181[183]^and_result181[184]^and_result181[185]^and_result181[186]^and_result181[187]^and_result181[188]^and_result181[189]^and_result181[190]^and_result181[191]^and_result181[192]^and_result181[193]^and_result181[194]^and_result181[195]^and_result181[196]^and_result181[197]^and_result181[198]^and_result181[199]^and_result181[200]^and_result181[201]^and_result181[202]^and_result181[203]^and_result181[204]^and_result181[205]^and_result181[206]^and_result181[207]^and_result181[208]^and_result181[209]^and_result181[210]^and_result181[211]^and_result181[212]^and_result181[213]^and_result181[214]^and_result181[215]^and_result181[216]^and_result181[217]^and_result181[218]^and_result181[219]^and_result181[220]^and_result181[221]^and_result181[222]^and_result181[223]^and_result181[224]^and_result181[225]^and_result181[226]^and_result181[227]^and_result181[228]^and_result181[229]^and_result181[230]^and_result181[231]^and_result181[232]^and_result181[233]^and_result181[234]^and_result181[235]^and_result181[236]^and_result181[237]^and_result181[238]^and_result181[239]^and_result181[240]^and_result181[241]^and_result181[242]^and_result181[243]^and_result181[244]^and_result181[245]^and_result181[246]^and_result181[247]^and_result181[248]^and_result181[249]^and_result181[250]^and_result181[251]^and_result181[252]^and_result181[253]^and_result181[254];
assign key[182]=and_result182[0]^and_result182[1]^and_result182[2]^and_result182[3]^and_result182[4]^and_result182[5]^and_result182[6]^and_result182[7]^and_result182[8]^and_result182[9]^and_result182[10]^and_result182[11]^and_result182[12]^and_result182[13]^and_result182[14]^and_result182[15]^and_result182[16]^and_result182[17]^and_result182[18]^and_result182[19]^and_result182[20]^and_result182[21]^and_result182[22]^and_result182[23]^and_result182[24]^and_result182[25]^and_result182[26]^and_result182[27]^and_result182[28]^and_result182[29]^and_result182[30]^and_result182[31]^and_result182[32]^and_result182[33]^and_result182[34]^and_result182[35]^and_result182[36]^and_result182[37]^and_result182[38]^and_result182[39]^and_result182[40]^and_result182[41]^and_result182[42]^and_result182[43]^and_result182[44]^and_result182[45]^and_result182[46]^and_result182[47]^and_result182[48]^and_result182[49]^and_result182[50]^and_result182[51]^and_result182[52]^and_result182[53]^and_result182[54]^and_result182[55]^and_result182[56]^and_result182[57]^and_result182[58]^and_result182[59]^and_result182[60]^and_result182[61]^and_result182[62]^and_result182[63]^and_result182[64]^and_result182[65]^and_result182[66]^and_result182[67]^and_result182[68]^and_result182[69]^and_result182[70]^and_result182[71]^and_result182[72]^and_result182[73]^and_result182[74]^and_result182[75]^and_result182[76]^and_result182[77]^and_result182[78]^and_result182[79]^and_result182[80]^and_result182[81]^and_result182[82]^and_result182[83]^and_result182[84]^and_result182[85]^and_result182[86]^and_result182[87]^and_result182[88]^and_result182[89]^and_result182[90]^and_result182[91]^and_result182[92]^and_result182[93]^and_result182[94]^and_result182[95]^and_result182[96]^and_result182[97]^and_result182[98]^and_result182[99]^and_result182[100]^and_result182[101]^and_result182[102]^and_result182[103]^and_result182[104]^and_result182[105]^and_result182[106]^and_result182[107]^and_result182[108]^and_result182[109]^and_result182[110]^and_result182[111]^and_result182[112]^and_result182[113]^and_result182[114]^and_result182[115]^and_result182[116]^and_result182[117]^and_result182[118]^and_result182[119]^and_result182[120]^and_result182[121]^and_result182[122]^and_result182[123]^and_result182[124]^and_result182[125]^and_result182[126]^and_result182[127]^and_result182[128]^and_result182[129]^and_result182[130]^and_result182[131]^and_result182[132]^and_result182[133]^and_result182[134]^and_result182[135]^and_result182[136]^and_result182[137]^and_result182[138]^and_result182[139]^and_result182[140]^and_result182[141]^and_result182[142]^and_result182[143]^and_result182[144]^and_result182[145]^and_result182[146]^and_result182[147]^and_result182[148]^and_result182[149]^and_result182[150]^and_result182[151]^and_result182[152]^and_result182[153]^and_result182[154]^and_result182[155]^and_result182[156]^and_result182[157]^and_result182[158]^and_result182[159]^and_result182[160]^and_result182[161]^and_result182[162]^and_result182[163]^and_result182[164]^and_result182[165]^and_result182[166]^and_result182[167]^and_result182[168]^and_result182[169]^and_result182[170]^and_result182[171]^and_result182[172]^and_result182[173]^and_result182[174]^and_result182[175]^and_result182[176]^and_result182[177]^and_result182[178]^and_result182[179]^and_result182[180]^and_result182[181]^and_result182[182]^and_result182[183]^and_result182[184]^and_result182[185]^and_result182[186]^and_result182[187]^and_result182[188]^and_result182[189]^and_result182[190]^and_result182[191]^and_result182[192]^and_result182[193]^and_result182[194]^and_result182[195]^and_result182[196]^and_result182[197]^and_result182[198]^and_result182[199]^and_result182[200]^and_result182[201]^and_result182[202]^and_result182[203]^and_result182[204]^and_result182[205]^and_result182[206]^and_result182[207]^and_result182[208]^and_result182[209]^and_result182[210]^and_result182[211]^and_result182[212]^and_result182[213]^and_result182[214]^and_result182[215]^and_result182[216]^and_result182[217]^and_result182[218]^and_result182[219]^and_result182[220]^and_result182[221]^and_result182[222]^and_result182[223]^and_result182[224]^and_result182[225]^and_result182[226]^and_result182[227]^and_result182[228]^and_result182[229]^and_result182[230]^and_result182[231]^and_result182[232]^and_result182[233]^and_result182[234]^and_result182[235]^and_result182[236]^and_result182[237]^and_result182[238]^and_result182[239]^and_result182[240]^and_result182[241]^and_result182[242]^and_result182[243]^and_result182[244]^and_result182[245]^and_result182[246]^and_result182[247]^and_result182[248]^and_result182[249]^and_result182[250]^and_result182[251]^and_result182[252]^and_result182[253]^and_result182[254];
assign key[183]=and_result183[0]^and_result183[1]^and_result183[2]^and_result183[3]^and_result183[4]^and_result183[5]^and_result183[6]^and_result183[7]^and_result183[8]^and_result183[9]^and_result183[10]^and_result183[11]^and_result183[12]^and_result183[13]^and_result183[14]^and_result183[15]^and_result183[16]^and_result183[17]^and_result183[18]^and_result183[19]^and_result183[20]^and_result183[21]^and_result183[22]^and_result183[23]^and_result183[24]^and_result183[25]^and_result183[26]^and_result183[27]^and_result183[28]^and_result183[29]^and_result183[30]^and_result183[31]^and_result183[32]^and_result183[33]^and_result183[34]^and_result183[35]^and_result183[36]^and_result183[37]^and_result183[38]^and_result183[39]^and_result183[40]^and_result183[41]^and_result183[42]^and_result183[43]^and_result183[44]^and_result183[45]^and_result183[46]^and_result183[47]^and_result183[48]^and_result183[49]^and_result183[50]^and_result183[51]^and_result183[52]^and_result183[53]^and_result183[54]^and_result183[55]^and_result183[56]^and_result183[57]^and_result183[58]^and_result183[59]^and_result183[60]^and_result183[61]^and_result183[62]^and_result183[63]^and_result183[64]^and_result183[65]^and_result183[66]^and_result183[67]^and_result183[68]^and_result183[69]^and_result183[70]^and_result183[71]^and_result183[72]^and_result183[73]^and_result183[74]^and_result183[75]^and_result183[76]^and_result183[77]^and_result183[78]^and_result183[79]^and_result183[80]^and_result183[81]^and_result183[82]^and_result183[83]^and_result183[84]^and_result183[85]^and_result183[86]^and_result183[87]^and_result183[88]^and_result183[89]^and_result183[90]^and_result183[91]^and_result183[92]^and_result183[93]^and_result183[94]^and_result183[95]^and_result183[96]^and_result183[97]^and_result183[98]^and_result183[99]^and_result183[100]^and_result183[101]^and_result183[102]^and_result183[103]^and_result183[104]^and_result183[105]^and_result183[106]^and_result183[107]^and_result183[108]^and_result183[109]^and_result183[110]^and_result183[111]^and_result183[112]^and_result183[113]^and_result183[114]^and_result183[115]^and_result183[116]^and_result183[117]^and_result183[118]^and_result183[119]^and_result183[120]^and_result183[121]^and_result183[122]^and_result183[123]^and_result183[124]^and_result183[125]^and_result183[126]^and_result183[127]^and_result183[128]^and_result183[129]^and_result183[130]^and_result183[131]^and_result183[132]^and_result183[133]^and_result183[134]^and_result183[135]^and_result183[136]^and_result183[137]^and_result183[138]^and_result183[139]^and_result183[140]^and_result183[141]^and_result183[142]^and_result183[143]^and_result183[144]^and_result183[145]^and_result183[146]^and_result183[147]^and_result183[148]^and_result183[149]^and_result183[150]^and_result183[151]^and_result183[152]^and_result183[153]^and_result183[154]^and_result183[155]^and_result183[156]^and_result183[157]^and_result183[158]^and_result183[159]^and_result183[160]^and_result183[161]^and_result183[162]^and_result183[163]^and_result183[164]^and_result183[165]^and_result183[166]^and_result183[167]^and_result183[168]^and_result183[169]^and_result183[170]^and_result183[171]^and_result183[172]^and_result183[173]^and_result183[174]^and_result183[175]^and_result183[176]^and_result183[177]^and_result183[178]^and_result183[179]^and_result183[180]^and_result183[181]^and_result183[182]^and_result183[183]^and_result183[184]^and_result183[185]^and_result183[186]^and_result183[187]^and_result183[188]^and_result183[189]^and_result183[190]^and_result183[191]^and_result183[192]^and_result183[193]^and_result183[194]^and_result183[195]^and_result183[196]^and_result183[197]^and_result183[198]^and_result183[199]^and_result183[200]^and_result183[201]^and_result183[202]^and_result183[203]^and_result183[204]^and_result183[205]^and_result183[206]^and_result183[207]^and_result183[208]^and_result183[209]^and_result183[210]^and_result183[211]^and_result183[212]^and_result183[213]^and_result183[214]^and_result183[215]^and_result183[216]^and_result183[217]^and_result183[218]^and_result183[219]^and_result183[220]^and_result183[221]^and_result183[222]^and_result183[223]^and_result183[224]^and_result183[225]^and_result183[226]^and_result183[227]^and_result183[228]^and_result183[229]^and_result183[230]^and_result183[231]^and_result183[232]^and_result183[233]^and_result183[234]^and_result183[235]^and_result183[236]^and_result183[237]^and_result183[238]^and_result183[239]^and_result183[240]^and_result183[241]^and_result183[242]^and_result183[243]^and_result183[244]^and_result183[245]^and_result183[246]^and_result183[247]^and_result183[248]^and_result183[249]^and_result183[250]^and_result183[251]^and_result183[252]^and_result183[253]^and_result183[254];
assign key[184]=and_result184[0]^and_result184[1]^and_result184[2]^and_result184[3]^and_result184[4]^and_result184[5]^and_result184[6]^and_result184[7]^and_result184[8]^and_result184[9]^and_result184[10]^and_result184[11]^and_result184[12]^and_result184[13]^and_result184[14]^and_result184[15]^and_result184[16]^and_result184[17]^and_result184[18]^and_result184[19]^and_result184[20]^and_result184[21]^and_result184[22]^and_result184[23]^and_result184[24]^and_result184[25]^and_result184[26]^and_result184[27]^and_result184[28]^and_result184[29]^and_result184[30]^and_result184[31]^and_result184[32]^and_result184[33]^and_result184[34]^and_result184[35]^and_result184[36]^and_result184[37]^and_result184[38]^and_result184[39]^and_result184[40]^and_result184[41]^and_result184[42]^and_result184[43]^and_result184[44]^and_result184[45]^and_result184[46]^and_result184[47]^and_result184[48]^and_result184[49]^and_result184[50]^and_result184[51]^and_result184[52]^and_result184[53]^and_result184[54]^and_result184[55]^and_result184[56]^and_result184[57]^and_result184[58]^and_result184[59]^and_result184[60]^and_result184[61]^and_result184[62]^and_result184[63]^and_result184[64]^and_result184[65]^and_result184[66]^and_result184[67]^and_result184[68]^and_result184[69]^and_result184[70]^and_result184[71]^and_result184[72]^and_result184[73]^and_result184[74]^and_result184[75]^and_result184[76]^and_result184[77]^and_result184[78]^and_result184[79]^and_result184[80]^and_result184[81]^and_result184[82]^and_result184[83]^and_result184[84]^and_result184[85]^and_result184[86]^and_result184[87]^and_result184[88]^and_result184[89]^and_result184[90]^and_result184[91]^and_result184[92]^and_result184[93]^and_result184[94]^and_result184[95]^and_result184[96]^and_result184[97]^and_result184[98]^and_result184[99]^and_result184[100]^and_result184[101]^and_result184[102]^and_result184[103]^and_result184[104]^and_result184[105]^and_result184[106]^and_result184[107]^and_result184[108]^and_result184[109]^and_result184[110]^and_result184[111]^and_result184[112]^and_result184[113]^and_result184[114]^and_result184[115]^and_result184[116]^and_result184[117]^and_result184[118]^and_result184[119]^and_result184[120]^and_result184[121]^and_result184[122]^and_result184[123]^and_result184[124]^and_result184[125]^and_result184[126]^and_result184[127]^and_result184[128]^and_result184[129]^and_result184[130]^and_result184[131]^and_result184[132]^and_result184[133]^and_result184[134]^and_result184[135]^and_result184[136]^and_result184[137]^and_result184[138]^and_result184[139]^and_result184[140]^and_result184[141]^and_result184[142]^and_result184[143]^and_result184[144]^and_result184[145]^and_result184[146]^and_result184[147]^and_result184[148]^and_result184[149]^and_result184[150]^and_result184[151]^and_result184[152]^and_result184[153]^and_result184[154]^and_result184[155]^and_result184[156]^and_result184[157]^and_result184[158]^and_result184[159]^and_result184[160]^and_result184[161]^and_result184[162]^and_result184[163]^and_result184[164]^and_result184[165]^and_result184[166]^and_result184[167]^and_result184[168]^and_result184[169]^and_result184[170]^and_result184[171]^and_result184[172]^and_result184[173]^and_result184[174]^and_result184[175]^and_result184[176]^and_result184[177]^and_result184[178]^and_result184[179]^and_result184[180]^and_result184[181]^and_result184[182]^and_result184[183]^and_result184[184]^and_result184[185]^and_result184[186]^and_result184[187]^and_result184[188]^and_result184[189]^and_result184[190]^and_result184[191]^and_result184[192]^and_result184[193]^and_result184[194]^and_result184[195]^and_result184[196]^and_result184[197]^and_result184[198]^and_result184[199]^and_result184[200]^and_result184[201]^and_result184[202]^and_result184[203]^and_result184[204]^and_result184[205]^and_result184[206]^and_result184[207]^and_result184[208]^and_result184[209]^and_result184[210]^and_result184[211]^and_result184[212]^and_result184[213]^and_result184[214]^and_result184[215]^and_result184[216]^and_result184[217]^and_result184[218]^and_result184[219]^and_result184[220]^and_result184[221]^and_result184[222]^and_result184[223]^and_result184[224]^and_result184[225]^and_result184[226]^and_result184[227]^and_result184[228]^and_result184[229]^and_result184[230]^and_result184[231]^and_result184[232]^and_result184[233]^and_result184[234]^and_result184[235]^and_result184[236]^and_result184[237]^and_result184[238]^and_result184[239]^and_result184[240]^and_result184[241]^and_result184[242]^and_result184[243]^and_result184[244]^and_result184[245]^and_result184[246]^and_result184[247]^and_result184[248]^and_result184[249]^and_result184[250]^and_result184[251]^and_result184[252]^and_result184[253]^and_result184[254];
assign key[185]=and_result185[0]^and_result185[1]^and_result185[2]^and_result185[3]^and_result185[4]^and_result185[5]^and_result185[6]^and_result185[7]^and_result185[8]^and_result185[9]^and_result185[10]^and_result185[11]^and_result185[12]^and_result185[13]^and_result185[14]^and_result185[15]^and_result185[16]^and_result185[17]^and_result185[18]^and_result185[19]^and_result185[20]^and_result185[21]^and_result185[22]^and_result185[23]^and_result185[24]^and_result185[25]^and_result185[26]^and_result185[27]^and_result185[28]^and_result185[29]^and_result185[30]^and_result185[31]^and_result185[32]^and_result185[33]^and_result185[34]^and_result185[35]^and_result185[36]^and_result185[37]^and_result185[38]^and_result185[39]^and_result185[40]^and_result185[41]^and_result185[42]^and_result185[43]^and_result185[44]^and_result185[45]^and_result185[46]^and_result185[47]^and_result185[48]^and_result185[49]^and_result185[50]^and_result185[51]^and_result185[52]^and_result185[53]^and_result185[54]^and_result185[55]^and_result185[56]^and_result185[57]^and_result185[58]^and_result185[59]^and_result185[60]^and_result185[61]^and_result185[62]^and_result185[63]^and_result185[64]^and_result185[65]^and_result185[66]^and_result185[67]^and_result185[68]^and_result185[69]^and_result185[70]^and_result185[71]^and_result185[72]^and_result185[73]^and_result185[74]^and_result185[75]^and_result185[76]^and_result185[77]^and_result185[78]^and_result185[79]^and_result185[80]^and_result185[81]^and_result185[82]^and_result185[83]^and_result185[84]^and_result185[85]^and_result185[86]^and_result185[87]^and_result185[88]^and_result185[89]^and_result185[90]^and_result185[91]^and_result185[92]^and_result185[93]^and_result185[94]^and_result185[95]^and_result185[96]^and_result185[97]^and_result185[98]^and_result185[99]^and_result185[100]^and_result185[101]^and_result185[102]^and_result185[103]^and_result185[104]^and_result185[105]^and_result185[106]^and_result185[107]^and_result185[108]^and_result185[109]^and_result185[110]^and_result185[111]^and_result185[112]^and_result185[113]^and_result185[114]^and_result185[115]^and_result185[116]^and_result185[117]^and_result185[118]^and_result185[119]^and_result185[120]^and_result185[121]^and_result185[122]^and_result185[123]^and_result185[124]^and_result185[125]^and_result185[126]^and_result185[127]^and_result185[128]^and_result185[129]^and_result185[130]^and_result185[131]^and_result185[132]^and_result185[133]^and_result185[134]^and_result185[135]^and_result185[136]^and_result185[137]^and_result185[138]^and_result185[139]^and_result185[140]^and_result185[141]^and_result185[142]^and_result185[143]^and_result185[144]^and_result185[145]^and_result185[146]^and_result185[147]^and_result185[148]^and_result185[149]^and_result185[150]^and_result185[151]^and_result185[152]^and_result185[153]^and_result185[154]^and_result185[155]^and_result185[156]^and_result185[157]^and_result185[158]^and_result185[159]^and_result185[160]^and_result185[161]^and_result185[162]^and_result185[163]^and_result185[164]^and_result185[165]^and_result185[166]^and_result185[167]^and_result185[168]^and_result185[169]^and_result185[170]^and_result185[171]^and_result185[172]^and_result185[173]^and_result185[174]^and_result185[175]^and_result185[176]^and_result185[177]^and_result185[178]^and_result185[179]^and_result185[180]^and_result185[181]^and_result185[182]^and_result185[183]^and_result185[184]^and_result185[185]^and_result185[186]^and_result185[187]^and_result185[188]^and_result185[189]^and_result185[190]^and_result185[191]^and_result185[192]^and_result185[193]^and_result185[194]^and_result185[195]^and_result185[196]^and_result185[197]^and_result185[198]^and_result185[199]^and_result185[200]^and_result185[201]^and_result185[202]^and_result185[203]^and_result185[204]^and_result185[205]^and_result185[206]^and_result185[207]^and_result185[208]^and_result185[209]^and_result185[210]^and_result185[211]^and_result185[212]^and_result185[213]^and_result185[214]^and_result185[215]^and_result185[216]^and_result185[217]^and_result185[218]^and_result185[219]^and_result185[220]^and_result185[221]^and_result185[222]^and_result185[223]^and_result185[224]^and_result185[225]^and_result185[226]^and_result185[227]^and_result185[228]^and_result185[229]^and_result185[230]^and_result185[231]^and_result185[232]^and_result185[233]^and_result185[234]^and_result185[235]^and_result185[236]^and_result185[237]^and_result185[238]^and_result185[239]^and_result185[240]^and_result185[241]^and_result185[242]^and_result185[243]^and_result185[244]^and_result185[245]^and_result185[246]^and_result185[247]^and_result185[248]^and_result185[249]^and_result185[250]^and_result185[251]^and_result185[252]^and_result185[253]^and_result185[254];
assign key[186]=and_result186[0]^and_result186[1]^and_result186[2]^and_result186[3]^and_result186[4]^and_result186[5]^and_result186[6]^and_result186[7]^and_result186[8]^and_result186[9]^and_result186[10]^and_result186[11]^and_result186[12]^and_result186[13]^and_result186[14]^and_result186[15]^and_result186[16]^and_result186[17]^and_result186[18]^and_result186[19]^and_result186[20]^and_result186[21]^and_result186[22]^and_result186[23]^and_result186[24]^and_result186[25]^and_result186[26]^and_result186[27]^and_result186[28]^and_result186[29]^and_result186[30]^and_result186[31]^and_result186[32]^and_result186[33]^and_result186[34]^and_result186[35]^and_result186[36]^and_result186[37]^and_result186[38]^and_result186[39]^and_result186[40]^and_result186[41]^and_result186[42]^and_result186[43]^and_result186[44]^and_result186[45]^and_result186[46]^and_result186[47]^and_result186[48]^and_result186[49]^and_result186[50]^and_result186[51]^and_result186[52]^and_result186[53]^and_result186[54]^and_result186[55]^and_result186[56]^and_result186[57]^and_result186[58]^and_result186[59]^and_result186[60]^and_result186[61]^and_result186[62]^and_result186[63]^and_result186[64]^and_result186[65]^and_result186[66]^and_result186[67]^and_result186[68]^and_result186[69]^and_result186[70]^and_result186[71]^and_result186[72]^and_result186[73]^and_result186[74]^and_result186[75]^and_result186[76]^and_result186[77]^and_result186[78]^and_result186[79]^and_result186[80]^and_result186[81]^and_result186[82]^and_result186[83]^and_result186[84]^and_result186[85]^and_result186[86]^and_result186[87]^and_result186[88]^and_result186[89]^and_result186[90]^and_result186[91]^and_result186[92]^and_result186[93]^and_result186[94]^and_result186[95]^and_result186[96]^and_result186[97]^and_result186[98]^and_result186[99]^and_result186[100]^and_result186[101]^and_result186[102]^and_result186[103]^and_result186[104]^and_result186[105]^and_result186[106]^and_result186[107]^and_result186[108]^and_result186[109]^and_result186[110]^and_result186[111]^and_result186[112]^and_result186[113]^and_result186[114]^and_result186[115]^and_result186[116]^and_result186[117]^and_result186[118]^and_result186[119]^and_result186[120]^and_result186[121]^and_result186[122]^and_result186[123]^and_result186[124]^and_result186[125]^and_result186[126]^and_result186[127]^and_result186[128]^and_result186[129]^and_result186[130]^and_result186[131]^and_result186[132]^and_result186[133]^and_result186[134]^and_result186[135]^and_result186[136]^and_result186[137]^and_result186[138]^and_result186[139]^and_result186[140]^and_result186[141]^and_result186[142]^and_result186[143]^and_result186[144]^and_result186[145]^and_result186[146]^and_result186[147]^and_result186[148]^and_result186[149]^and_result186[150]^and_result186[151]^and_result186[152]^and_result186[153]^and_result186[154]^and_result186[155]^and_result186[156]^and_result186[157]^and_result186[158]^and_result186[159]^and_result186[160]^and_result186[161]^and_result186[162]^and_result186[163]^and_result186[164]^and_result186[165]^and_result186[166]^and_result186[167]^and_result186[168]^and_result186[169]^and_result186[170]^and_result186[171]^and_result186[172]^and_result186[173]^and_result186[174]^and_result186[175]^and_result186[176]^and_result186[177]^and_result186[178]^and_result186[179]^and_result186[180]^and_result186[181]^and_result186[182]^and_result186[183]^and_result186[184]^and_result186[185]^and_result186[186]^and_result186[187]^and_result186[188]^and_result186[189]^and_result186[190]^and_result186[191]^and_result186[192]^and_result186[193]^and_result186[194]^and_result186[195]^and_result186[196]^and_result186[197]^and_result186[198]^and_result186[199]^and_result186[200]^and_result186[201]^and_result186[202]^and_result186[203]^and_result186[204]^and_result186[205]^and_result186[206]^and_result186[207]^and_result186[208]^and_result186[209]^and_result186[210]^and_result186[211]^and_result186[212]^and_result186[213]^and_result186[214]^and_result186[215]^and_result186[216]^and_result186[217]^and_result186[218]^and_result186[219]^and_result186[220]^and_result186[221]^and_result186[222]^and_result186[223]^and_result186[224]^and_result186[225]^and_result186[226]^and_result186[227]^and_result186[228]^and_result186[229]^and_result186[230]^and_result186[231]^and_result186[232]^and_result186[233]^and_result186[234]^and_result186[235]^and_result186[236]^and_result186[237]^and_result186[238]^and_result186[239]^and_result186[240]^and_result186[241]^and_result186[242]^and_result186[243]^and_result186[244]^and_result186[245]^and_result186[246]^and_result186[247]^and_result186[248]^and_result186[249]^and_result186[250]^and_result186[251]^and_result186[252]^and_result186[253]^and_result186[254];
assign key[187]=and_result187[0]^and_result187[1]^and_result187[2]^and_result187[3]^and_result187[4]^and_result187[5]^and_result187[6]^and_result187[7]^and_result187[8]^and_result187[9]^and_result187[10]^and_result187[11]^and_result187[12]^and_result187[13]^and_result187[14]^and_result187[15]^and_result187[16]^and_result187[17]^and_result187[18]^and_result187[19]^and_result187[20]^and_result187[21]^and_result187[22]^and_result187[23]^and_result187[24]^and_result187[25]^and_result187[26]^and_result187[27]^and_result187[28]^and_result187[29]^and_result187[30]^and_result187[31]^and_result187[32]^and_result187[33]^and_result187[34]^and_result187[35]^and_result187[36]^and_result187[37]^and_result187[38]^and_result187[39]^and_result187[40]^and_result187[41]^and_result187[42]^and_result187[43]^and_result187[44]^and_result187[45]^and_result187[46]^and_result187[47]^and_result187[48]^and_result187[49]^and_result187[50]^and_result187[51]^and_result187[52]^and_result187[53]^and_result187[54]^and_result187[55]^and_result187[56]^and_result187[57]^and_result187[58]^and_result187[59]^and_result187[60]^and_result187[61]^and_result187[62]^and_result187[63]^and_result187[64]^and_result187[65]^and_result187[66]^and_result187[67]^and_result187[68]^and_result187[69]^and_result187[70]^and_result187[71]^and_result187[72]^and_result187[73]^and_result187[74]^and_result187[75]^and_result187[76]^and_result187[77]^and_result187[78]^and_result187[79]^and_result187[80]^and_result187[81]^and_result187[82]^and_result187[83]^and_result187[84]^and_result187[85]^and_result187[86]^and_result187[87]^and_result187[88]^and_result187[89]^and_result187[90]^and_result187[91]^and_result187[92]^and_result187[93]^and_result187[94]^and_result187[95]^and_result187[96]^and_result187[97]^and_result187[98]^and_result187[99]^and_result187[100]^and_result187[101]^and_result187[102]^and_result187[103]^and_result187[104]^and_result187[105]^and_result187[106]^and_result187[107]^and_result187[108]^and_result187[109]^and_result187[110]^and_result187[111]^and_result187[112]^and_result187[113]^and_result187[114]^and_result187[115]^and_result187[116]^and_result187[117]^and_result187[118]^and_result187[119]^and_result187[120]^and_result187[121]^and_result187[122]^and_result187[123]^and_result187[124]^and_result187[125]^and_result187[126]^and_result187[127]^and_result187[128]^and_result187[129]^and_result187[130]^and_result187[131]^and_result187[132]^and_result187[133]^and_result187[134]^and_result187[135]^and_result187[136]^and_result187[137]^and_result187[138]^and_result187[139]^and_result187[140]^and_result187[141]^and_result187[142]^and_result187[143]^and_result187[144]^and_result187[145]^and_result187[146]^and_result187[147]^and_result187[148]^and_result187[149]^and_result187[150]^and_result187[151]^and_result187[152]^and_result187[153]^and_result187[154]^and_result187[155]^and_result187[156]^and_result187[157]^and_result187[158]^and_result187[159]^and_result187[160]^and_result187[161]^and_result187[162]^and_result187[163]^and_result187[164]^and_result187[165]^and_result187[166]^and_result187[167]^and_result187[168]^and_result187[169]^and_result187[170]^and_result187[171]^and_result187[172]^and_result187[173]^and_result187[174]^and_result187[175]^and_result187[176]^and_result187[177]^and_result187[178]^and_result187[179]^and_result187[180]^and_result187[181]^and_result187[182]^and_result187[183]^and_result187[184]^and_result187[185]^and_result187[186]^and_result187[187]^and_result187[188]^and_result187[189]^and_result187[190]^and_result187[191]^and_result187[192]^and_result187[193]^and_result187[194]^and_result187[195]^and_result187[196]^and_result187[197]^and_result187[198]^and_result187[199]^and_result187[200]^and_result187[201]^and_result187[202]^and_result187[203]^and_result187[204]^and_result187[205]^and_result187[206]^and_result187[207]^and_result187[208]^and_result187[209]^and_result187[210]^and_result187[211]^and_result187[212]^and_result187[213]^and_result187[214]^and_result187[215]^and_result187[216]^and_result187[217]^and_result187[218]^and_result187[219]^and_result187[220]^and_result187[221]^and_result187[222]^and_result187[223]^and_result187[224]^and_result187[225]^and_result187[226]^and_result187[227]^and_result187[228]^and_result187[229]^and_result187[230]^and_result187[231]^and_result187[232]^and_result187[233]^and_result187[234]^and_result187[235]^and_result187[236]^and_result187[237]^and_result187[238]^and_result187[239]^and_result187[240]^and_result187[241]^and_result187[242]^and_result187[243]^and_result187[244]^and_result187[245]^and_result187[246]^and_result187[247]^and_result187[248]^and_result187[249]^and_result187[250]^and_result187[251]^and_result187[252]^and_result187[253]^and_result187[254];
assign key[188]=and_result188[0]^and_result188[1]^and_result188[2]^and_result188[3]^and_result188[4]^and_result188[5]^and_result188[6]^and_result188[7]^and_result188[8]^and_result188[9]^and_result188[10]^and_result188[11]^and_result188[12]^and_result188[13]^and_result188[14]^and_result188[15]^and_result188[16]^and_result188[17]^and_result188[18]^and_result188[19]^and_result188[20]^and_result188[21]^and_result188[22]^and_result188[23]^and_result188[24]^and_result188[25]^and_result188[26]^and_result188[27]^and_result188[28]^and_result188[29]^and_result188[30]^and_result188[31]^and_result188[32]^and_result188[33]^and_result188[34]^and_result188[35]^and_result188[36]^and_result188[37]^and_result188[38]^and_result188[39]^and_result188[40]^and_result188[41]^and_result188[42]^and_result188[43]^and_result188[44]^and_result188[45]^and_result188[46]^and_result188[47]^and_result188[48]^and_result188[49]^and_result188[50]^and_result188[51]^and_result188[52]^and_result188[53]^and_result188[54]^and_result188[55]^and_result188[56]^and_result188[57]^and_result188[58]^and_result188[59]^and_result188[60]^and_result188[61]^and_result188[62]^and_result188[63]^and_result188[64]^and_result188[65]^and_result188[66]^and_result188[67]^and_result188[68]^and_result188[69]^and_result188[70]^and_result188[71]^and_result188[72]^and_result188[73]^and_result188[74]^and_result188[75]^and_result188[76]^and_result188[77]^and_result188[78]^and_result188[79]^and_result188[80]^and_result188[81]^and_result188[82]^and_result188[83]^and_result188[84]^and_result188[85]^and_result188[86]^and_result188[87]^and_result188[88]^and_result188[89]^and_result188[90]^and_result188[91]^and_result188[92]^and_result188[93]^and_result188[94]^and_result188[95]^and_result188[96]^and_result188[97]^and_result188[98]^and_result188[99]^and_result188[100]^and_result188[101]^and_result188[102]^and_result188[103]^and_result188[104]^and_result188[105]^and_result188[106]^and_result188[107]^and_result188[108]^and_result188[109]^and_result188[110]^and_result188[111]^and_result188[112]^and_result188[113]^and_result188[114]^and_result188[115]^and_result188[116]^and_result188[117]^and_result188[118]^and_result188[119]^and_result188[120]^and_result188[121]^and_result188[122]^and_result188[123]^and_result188[124]^and_result188[125]^and_result188[126]^and_result188[127]^and_result188[128]^and_result188[129]^and_result188[130]^and_result188[131]^and_result188[132]^and_result188[133]^and_result188[134]^and_result188[135]^and_result188[136]^and_result188[137]^and_result188[138]^and_result188[139]^and_result188[140]^and_result188[141]^and_result188[142]^and_result188[143]^and_result188[144]^and_result188[145]^and_result188[146]^and_result188[147]^and_result188[148]^and_result188[149]^and_result188[150]^and_result188[151]^and_result188[152]^and_result188[153]^and_result188[154]^and_result188[155]^and_result188[156]^and_result188[157]^and_result188[158]^and_result188[159]^and_result188[160]^and_result188[161]^and_result188[162]^and_result188[163]^and_result188[164]^and_result188[165]^and_result188[166]^and_result188[167]^and_result188[168]^and_result188[169]^and_result188[170]^and_result188[171]^and_result188[172]^and_result188[173]^and_result188[174]^and_result188[175]^and_result188[176]^and_result188[177]^and_result188[178]^and_result188[179]^and_result188[180]^and_result188[181]^and_result188[182]^and_result188[183]^and_result188[184]^and_result188[185]^and_result188[186]^and_result188[187]^and_result188[188]^and_result188[189]^and_result188[190]^and_result188[191]^and_result188[192]^and_result188[193]^and_result188[194]^and_result188[195]^and_result188[196]^and_result188[197]^and_result188[198]^and_result188[199]^and_result188[200]^and_result188[201]^and_result188[202]^and_result188[203]^and_result188[204]^and_result188[205]^and_result188[206]^and_result188[207]^and_result188[208]^and_result188[209]^and_result188[210]^and_result188[211]^and_result188[212]^and_result188[213]^and_result188[214]^and_result188[215]^and_result188[216]^and_result188[217]^and_result188[218]^and_result188[219]^and_result188[220]^and_result188[221]^and_result188[222]^and_result188[223]^and_result188[224]^and_result188[225]^and_result188[226]^and_result188[227]^and_result188[228]^and_result188[229]^and_result188[230]^and_result188[231]^and_result188[232]^and_result188[233]^and_result188[234]^and_result188[235]^and_result188[236]^and_result188[237]^and_result188[238]^and_result188[239]^and_result188[240]^and_result188[241]^and_result188[242]^and_result188[243]^and_result188[244]^and_result188[245]^and_result188[246]^and_result188[247]^and_result188[248]^and_result188[249]^and_result188[250]^and_result188[251]^and_result188[252]^and_result188[253]^and_result188[254];
assign key[189]=and_result189[0]^and_result189[1]^and_result189[2]^and_result189[3]^and_result189[4]^and_result189[5]^and_result189[6]^and_result189[7]^and_result189[8]^and_result189[9]^and_result189[10]^and_result189[11]^and_result189[12]^and_result189[13]^and_result189[14]^and_result189[15]^and_result189[16]^and_result189[17]^and_result189[18]^and_result189[19]^and_result189[20]^and_result189[21]^and_result189[22]^and_result189[23]^and_result189[24]^and_result189[25]^and_result189[26]^and_result189[27]^and_result189[28]^and_result189[29]^and_result189[30]^and_result189[31]^and_result189[32]^and_result189[33]^and_result189[34]^and_result189[35]^and_result189[36]^and_result189[37]^and_result189[38]^and_result189[39]^and_result189[40]^and_result189[41]^and_result189[42]^and_result189[43]^and_result189[44]^and_result189[45]^and_result189[46]^and_result189[47]^and_result189[48]^and_result189[49]^and_result189[50]^and_result189[51]^and_result189[52]^and_result189[53]^and_result189[54]^and_result189[55]^and_result189[56]^and_result189[57]^and_result189[58]^and_result189[59]^and_result189[60]^and_result189[61]^and_result189[62]^and_result189[63]^and_result189[64]^and_result189[65]^and_result189[66]^and_result189[67]^and_result189[68]^and_result189[69]^and_result189[70]^and_result189[71]^and_result189[72]^and_result189[73]^and_result189[74]^and_result189[75]^and_result189[76]^and_result189[77]^and_result189[78]^and_result189[79]^and_result189[80]^and_result189[81]^and_result189[82]^and_result189[83]^and_result189[84]^and_result189[85]^and_result189[86]^and_result189[87]^and_result189[88]^and_result189[89]^and_result189[90]^and_result189[91]^and_result189[92]^and_result189[93]^and_result189[94]^and_result189[95]^and_result189[96]^and_result189[97]^and_result189[98]^and_result189[99]^and_result189[100]^and_result189[101]^and_result189[102]^and_result189[103]^and_result189[104]^and_result189[105]^and_result189[106]^and_result189[107]^and_result189[108]^and_result189[109]^and_result189[110]^and_result189[111]^and_result189[112]^and_result189[113]^and_result189[114]^and_result189[115]^and_result189[116]^and_result189[117]^and_result189[118]^and_result189[119]^and_result189[120]^and_result189[121]^and_result189[122]^and_result189[123]^and_result189[124]^and_result189[125]^and_result189[126]^and_result189[127]^and_result189[128]^and_result189[129]^and_result189[130]^and_result189[131]^and_result189[132]^and_result189[133]^and_result189[134]^and_result189[135]^and_result189[136]^and_result189[137]^and_result189[138]^and_result189[139]^and_result189[140]^and_result189[141]^and_result189[142]^and_result189[143]^and_result189[144]^and_result189[145]^and_result189[146]^and_result189[147]^and_result189[148]^and_result189[149]^and_result189[150]^and_result189[151]^and_result189[152]^and_result189[153]^and_result189[154]^and_result189[155]^and_result189[156]^and_result189[157]^and_result189[158]^and_result189[159]^and_result189[160]^and_result189[161]^and_result189[162]^and_result189[163]^and_result189[164]^and_result189[165]^and_result189[166]^and_result189[167]^and_result189[168]^and_result189[169]^and_result189[170]^and_result189[171]^and_result189[172]^and_result189[173]^and_result189[174]^and_result189[175]^and_result189[176]^and_result189[177]^and_result189[178]^and_result189[179]^and_result189[180]^and_result189[181]^and_result189[182]^and_result189[183]^and_result189[184]^and_result189[185]^and_result189[186]^and_result189[187]^and_result189[188]^and_result189[189]^and_result189[190]^and_result189[191]^and_result189[192]^and_result189[193]^and_result189[194]^and_result189[195]^and_result189[196]^and_result189[197]^and_result189[198]^and_result189[199]^and_result189[200]^and_result189[201]^and_result189[202]^and_result189[203]^and_result189[204]^and_result189[205]^and_result189[206]^and_result189[207]^and_result189[208]^and_result189[209]^and_result189[210]^and_result189[211]^and_result189[212]^and_result189[213]^and_result189[214]^and_result189[215]^and_result189[216]^and_result189[217]^and_result189[218]^and_result189[219]^and_result189[220]^and_result189[221]^and_result189[222]^and_result189[223]^and_result189[224]^and_result189[225]^and_result189[226]^and_result189[227]^and_result189[228]^and_result189[229]^and_result189[230]^and_result189[231]^and_result189[232]^and_result189[233]^and_result189[234]^and_result189[235]^and_result189[236]^and_result189[237]^and_result189[238]^and_result189[239]^and_result189[240]^and_result189[241]^and_result189[242]^and_result189[243]^and_result189[244]^and_result189[245]^and_result189[246]^and_result189[247]^and_result189[248]^and_result189[249]^and_result189[250]^and_result189[251]^and_result189[252]^and_result189[253]^and_result189[254];
assign key[190]=and_result190[0]^and_result190[1]^and_result190[2]^and_result190[3]^and_result190[4]^and_result190[5]^and_result190[6]^and_result190[7]^and_result190[8]^and_result190[9]^and_result190[10]^and_result190[11]^and_result190[12]^and_result190[13]^and_result190[14]^and_result190[15]^and_result190[16]^and_result190[17]^and_result190[18]^and_result190[19]^and_result190[20]^and_result190[21]^and_result190[22]^and_result190[23]^and_result190[24]^and_result190[25]^and_result190[26]^and_result190[27]^and_result190[28]^and_result190[29]^and_result190[30]^and_result190[31]^and_result190[32]^and_result190[33]^and_result190[34]^and_result190[35]^and_result190[36]^and_result190[37]^and_result190[38]^and_result190[39]^and_result190[40]^and_result190[41]^and_result190[42]^and_result190[43]^and_result190[44]^and_result190[45]^and_result190[46]^and_result190[47]^and_result190[48]^and_result190[49]^and_result190[50]^and_result190[51]^and_result190[52]^and_result190[53]^and_result190[54]^and_result190[55]^and_result190[56]^and_result190[57]^and_result190[58]^and_result190[59]^and_result190[60]^and_result190[61]^and_result190[62]^and_result190[63]^and_result190[64]^and_result190[65]^and_result190[66]^and_result190[67]^and_result190[68]^and_result190[69]^and_result190[70]^and_result190[71]^and_result190[72]^and_result190[73]^and_result190[74]^and_result190[75]^and_result190[76]^and_result190[77]^and_result190[78]^and_result190[79]^and_result190[80]^and_result190[81]^and_result190[82]^and_result190[83]^and_result190[84]^and_result190[85]^and_result190[86]^and_result190[87]^and_result190[88]^and_result190[89]^and_result190[90]^and_result190[91]^and_result190[92]^and_result190[93]^and_result190[94]^and_result190[95]^and_result190[96]^and_result190[97]^and_result190[98]^and_result190[99]^and_result190[100]^and_result190[101]^and_result190[102]^and_result190[103]^and_result190[104]^and_result190[105]^and_result190[106]^and_result190[107]^and_result190[108]^and_result190[109]^and_result190[110]^and_result190[111]^and_result190[112]^and_result190[113]^and_result190[114]^and_result190[115]^and_result190[116]^and_result190[117]^and_result190[118]^and_result190[119]^and_result190[120]^and_result190[121]^and_result190[122]^and_result190[123]^and_result190[124]^and_result190[125]^and_result190[126]^and_result190[127]^and_result190[128]^and_result190[129]^and_result190[130]^and_result190[131]^and_result190[132]^and_result190[133]^and_result190[134]^and_result190[135]^and_result190[136]^and_result190[137]^and_result190[138]^and_result190[139]^and_result190[140]^and_result190[141]^and_result190[142]^and_result190[143]^and_result190[144]^and_result190[145]^and_result190[146]^and_result190[147]^and_result190[148]^and_result190[149]^and_result190[150]^and_result190[151]^and_result190[152]^and_result190[153]^and_result190[154]^and_result190[155]^and_result190[156]^and_result190[157]^and_result190[158]^and_result190[159]^and_result190[160]^and_result190[161]^and_result190[162]^and_result190[163]^and_result190[164]^and_result190[165]^and_result190[166]^and_result190[167]^and_result190[168]^and_result190[169]^and_result190[170]^and_result190[171]^and_result190[172]^and_result190[173]^and_result190[174]^and_result190[175]^and_result190[176]^and_result190[177]^and_result190[178]^and_result190[179]^and_result190[180]^and_result190[181]^and_result190[182]^and_result190[183]^and_result190[184]^and_result190[185]^and_result190[186]^and_result190[187]^and_result190[188]^and_result190[189]^and_result190[190]^and_result190[191]^and_result190[192]^and_result190[193]^and_result190[194]^and_result190[195]^and_result190[196]^and_result190[197]^and_result190[198]^and_result190[199]^and_result190[200]^and_result190[201]^and_result190[202]^and_result190[203]^and_result190[204]^and_result190[205]^and_result190[206]^and_result190[207]^and_result190[208]^and_result190[209]^and_result190[210]^and_result190[211]^and_result190[212]^and_result190[213]^and_result190[214]^and_result190[215]^and_result190[216]^and_result190[217]^and_result190[218]^and_result190[219]^and_result190[220]^and_result190[221]^and_result190[222]^and_result190[223]^and_result190[224]^and_result190[225]^and_result190[226]^and_result190[227]^and_result190[228]^and_result190[229]^and_result190[230]^and_result190[231]^and_result190[232]^and_result190[233]^and_result190[234]^and_result190[235]^and_result190[236]^and_result190[237]^and_result190[238]^and_result190[239]^and_result190[240]^and_result190[241]^and_result190[242]^and_result190[243]^and_result190[244]^and_result190[245]^and_result190[246]^and_result190[247]^and_result190[248]^and_result190[249]^and_result190[250]^and_result190[251]^and_result190[252]^and_result190[253]^and_result190[254];
assign key[191]=and_result191[0]^and_result191[1]^and_result191[2]^and_result191[3]^and_result191[4]^and_result191[5]^and_result191[6]^and_result191[7]^and_result191[8]^and_result191[9]^and_result191[10]^and_result191[11]^and_result191[12]^and_result191[13]^and_result191[14]^and_result191[15]^and_result191[16]^and_result191[17]^and_result191[18]^and_result191[19]^and_result191[20]^and_result191[21]^and_result191[22]^and_result191[23]^and_result191[24]^and_result191[25]^and_result191[26]^and_result191[27]^and_result191[28]^and_result191[29]^and_result191[30]^and_result191[31]^and_result191[32]^and_result191[33]^and_result191[34]^and_result191[35]^and_result191[36]^and_result191[37]^and_result191[38]^and_result191[39]^and_result191[40]^and_result191[41]^and_result191[42]^and_result191[43]^and_result191[44]^and_result191[45]^and_result191[46]^and_result191[47]^and_result191[48]^and_result191[49]^and_result191[50]^and_result191[51]^and_result191[52]^and_result191[53]^and_result191[54]^and_result191[55]^and_result191[56]^and_result191[57]^and_result191[58]^and_result191[59]^and_result191[60]^and_result191[61]^and_result191[62]^and_result191[63]^and_result191[64]^and_result191[65]^and_result191[66]^and_result191[67]^and_result191[68]^and_result191[69]^and_result191[70]^and_result191[71]^and_result191[72]^and_result191[73]^and_result191[74]^and_result191[75]^and_result191[76]^and_result191[77]^and_result191[78]^and_result191[79]^and_result191[80]^and_result191[81]^and_result191[82]^and_result191[83]^and_result191[84]^and_result191[85]^and_result191[86]^and_result191[87]^and_result191[88]^and_result191[89]^and_result191[90]^and_result191[91]^and_result191[92]^and_result191[93]^and_result191[94]^and_result191[95]^and_result191[96]^and_result191[97]^and_result191[98]^and_result191[99]^and_result191[100]^and_result191[101]^and_result191[102]^and_result191[103]^and_result191[104]^and_result191[105]^and_result191[106]^and_result191[107]^and_result191[108]^and_result191[109]^and_result191[110]^and_result191[111]^and_result191[112]^and_result191[113]^and_result191[114]^and_result191[115]^and_result191[116]^and_result191[117]^and_result191[118]^and_result191[119]^and_result191[120]^and_result191[121]^and_result191[122]^and_result191[123]^and_result191[124]^and_result191[125]^and_result191[126]^and_result191[127]^and_result191[128]^and_result191[129]^and_result191[130]^and_result191[131]^and_result191[132]^and_result191[133]^and_result191[134]^and_result191[135]^and_result191[136]^and_result191[137]^and_result191[138]^and_result191[139]^and_result191[140]^and_result191[141]^and_result191[142]^and_result191[143]^and_result191[144]^and_result191[145]^and_result191[146]^and_result191[147]^and_result191[148]^and_result191[149]^and_result191[150]^and_result191[151]^and_result191[152]^and_result191[153]^and_result191[154]^and_result191[155]^and_result191[156]^and_result191[157]^and_result191[158]^and_result191[159]^and_result191[160]^and_result191[161]^and_result191[162]^and_result191[163]^and_result191[164]^and_result191[165]^and_result191[166]^and_result191[167]^and_result191[168]^and_result191[169]^and_result191[170]^and_result191[171]^and_result191[172]^and_result191[173]^and_result191[174]^and_result191[175]^and_result191[176]^and_result191[177]^and_result191[178]^and_result191[179]^and_result191[180]^and_result191[181]^and_result191[182]^and_result191[183]^and_result191[184]^and_result191[185]^and_result191[186]^and_result191[187]^and_result191[188]^and_result191[189]^and_result191[190]^and_result191[191]^and_result191[192]^and_result191[193]^and_result191[194]^and_result191[195]^and_result191[196]^and_result191[197]^and_result191[198]^and_result191[199]^and_result191[200]^and_result191[201]^and_result191[202]^and_result191[203]^and_result191[204]^and_result191[205]^and_result191[206]^and_result191[207]^and_result191[208]^and_result191[209]^and_result191[210]^and_result191[211]^and_result191[212]^and_result191[213]^and_result191[214]^and_result191[215]^and_result191[216]^and_result191[217]^and_result191[218]^and_result191[219]^and_result191[220]^and_result191[221]^and_result191[222]^and_result191[223]^and_result191[224]^and_result191[225]^and_result191[226]^and_result191[227]^and_result191[228]^and_result191[229]^and_result191[230]^and_result191[231]^and_result191[232]^and_result191[233]^and_result191[234]^and_result191[235]^and_result191[236]^and_result191[237]^and_result191[238]^and_result191[239]^and_result191[240]^and_result191[241]^and_result191[242]^and_result191[243]^and_result191[244]^and_result191[245]^and_result191[246]^and_result191[247]^and_result191[248]^and_result191[249]^and_result191[250]^and_result191[251]^and_result191[252]^and_result191[253]^and_result191[254];
assign key[192]=and_result192[0]^and_result192[1]^and_result192[2]^and_result192[3]^and_result192[4]^and_result192[5]^and_result192[6]^and_result192[7]^and_result192[8]^and_result192[9]^and_result192[10]^and_result192[11]^and_result192[12]^and_result192[13]^and_result192[14]^and_result192[15]^and_result192[16]^and_result192[17]^and_result192[18]^and_result192[19]^and_result192[20]^and_result192[21]^and_result192[22]^and_result192[23]^and_result192[24]^and_result192[25]^and_result192[26]^and_result192[27]^and_result192[28]^and_result192[29]^and_result192[30]^and_result192[31]^and_result192[32]^and_result192[33]^and_result192[34]^and_result192[35]^and_result192[36]^and_result192[37]^and_result192[38]^and_result192[39]^and_result192[40]^and_result192[41]^and_result192[42]^and_result192[43]^and_result192[44]^and_result192[45]^and_result192[46]^and_result192[47]^and_result192[48]^and_result192[49]^and_result192[50]^and_result192[51]^and_result192[52]^and_result192[53]^and_result192[54]^and_result192[55]^and_result192[56]^and_result192[57]^and_result192[58]^and_result192[59]^and_result192[60]^and_result192[61]^and_result192[62]^and_result192[63]^and_result192[64]^and_result192[65]^and_result192[66]^and_result192[67]^and_result192[68]^and_result192[69]^and_result192[70]^and_result192[71]^and_result192[72]^and_result192[73]^and_result192[74]^and_result192[75]^and_result192[76]^and_result192[77]^and_result192[78]^and_result192[79]^and_result192[80]^and_result192[81]^and_result192[82]^and_result192[83]^and_result192[84]^and_result192[85]^and_result192[86]^and_result192[87]^and_result192[88]^and_result192[89]^and_result192[90]^and_result192[91]^and_result192[92]^and_result192[93]^and_result192[94]^and_result192[95]^and_result192[96]^and_result192[97]^and_result192[98]^and_result192[99]^and_result192[100]^and_result192[101]^and_result192[102]^and_result192[103]^and_result192[104]^and_result192[105]^and_result192[106]^and_result192[107]^and_result192[108]^and_result192[109]^and_result192[110]^and_result192[111]^and_result192[112]^and_result192[113]^and_result192[114]^and_result192[115]^and_result192[116]^and_result192[117]^and_result192[118]^and_result192[119]^and_result192[120]^and_result192[121]^and_result192[122]^and_result192[123]^and_result192[124]^and_result192[125]^and_result192[126]^and_result192[127]^and_result192[128]^and_result192[129]^and_result192[130]^and_result192[131]^and_result192[132]^and_result192[133]^and_result192[134]^and_result192[135]^and_result192[136]^and_result192[137]^and_result192[138]^and_result192[139]^and_result192[140]^and_result192[141]^and_result192[142]^and_result192[143]^and_result192[144]^and_result192[145]^and_result192[146]^and_result192[147]^and_result192[148]^and_result192[149]^and_result192[150]^and_result192[151]^and_result192[152]^and_result192[153]^and_result192[154]^and_result192[155]^and_result192[156]^and_result192[157]^and_result192[158]^and_result192[159]^and_result192[160]^and_result192[161]^and_result192[162]^and_result192[163]^and_result192[164]^and_result192[165]^and_result192[166]^and_result192[167]^and_result192[168]^and_result192[169]^and_result192[170]^and_result192[171]^and_result192[172]^and_result192[173]^and_result192[174]^and_result192[175]^and_result192[176]^and_result192[177]^and_result192[178]^and_result192[179]^and_result192[180]^and_result192[181]^and_result192[182]^and_result192[183]^and_result192[184]^and_result192[185]^and_result192[186]^and_result192[187]^and_result192[188]^and_result192[189]^and_result192[190]^and_result192[191]^and_result192[192]^and_result192[193]^and_result192[194]^and_result192[195]^and_result192[196]^and_result192[197]^and_result192[198]^and_result192[199]^and_result192[200]^and_result192[201]^and_result192[202]^and_result192[203]^and_result192[204]^and_result192[205]^and_result192[206]^and_result192[207]^and_result192[208]^and_result192[209]^and_result192[210]^and_result192[211]^and_result192[212]^and_result192[213]^and_result192[214]^and_result192[215]^and_result192[216]^and_result192[217]^and_result192[218]^and_result192[219]^and_result192[220]^and_result192[221]^and_result192[222]^and_result192[223]^and_result192[224]^and_result192[225]^and_result192[226]^and_result192[227]^and_result192[228]^and_result192[229]^and_result192[230]^and_result192[231]^and_result192[232]^and_result192[233]^and_result192[234]^and_result192[235]^and_result192[236]^and_result192[237]^and_result192[238]^and_result192[239]^and_result192[240]^and_result192[241]^and_result192[242]^and_result192[243]^and_result192[244]^and_result192[245]^and_result192[246]^and_result192[247]^and_result192[248]^and_result192[249]^and_result192[250]^and_result192[251]^and_result192[252]^and_result192[253]^and_result192[254];
assign key[193]=and_result193[0]^and_result193[1]^and_result193[2]^and_result193[3]^and_result193[4]^and_result193[5]^and_result193[6]^and_result193[7]^and_result193[8]^and_result193[9]^and_result193[10]^and_result193[11]^and_result193[12]^and_result193[13]^and_result193[14]^and_result193[15]^and_result193[16]^and_result193[17]^and_result193[18]^and_result193[19]^and_result193[20]^and_result193[21]^and_result193[22]^and_result193[23]^and_result193[24]^and_result193[25]^and_result193[26]^and_result193[27]^and_result193[28]^and_result193[29]^and_result193[30]^and_result193[31]^and_result193[32]^and_result193[33]^and_result193[34]^and_result193[35]^and_result193[36]^and_result193[37]^and_result193[38]^and_result193[39]^and_result193[40]^and_result193[41]^and_result193[42]^and_result193[43]^and_result193[44]^and_result193[45]^and_result193[46]^and_result193[47]^and_result193[48]^and_result193[49]^and_result193[50]^and_result193[51]^and_result193[52]^and_result193[53]^and_result193[54]^and_result193[55]^and_result193[56]^and_result193[57]^and_result193[58]^and_result193[59]^and_result193[60]^and_result193[61]^and_result193[62]^and_result193[63]^and_result193[64]^and_result193[65]^and_result193[66]^and_result193[67]^and_result193[68]^and_result193[69]^and_result193[70]^and_result193[71]^and_result193[72]^and_result193[73]^and_result193[74]^and_result193[75]^and_result193[76]^and_result193[77]^and_result193[78]^and_result193[79]^and_result193[80]^and_result193[81]^and_result193[82]^and_result193[83]^and_result193[84]^and_result193[85]^and_result193[86]^and_result193[87]^and_result193[88]^and_result193[89]^and_result193[90]^and_result193[91]^and_result193[92]^and_result193[93]^and_result193[94]^and_result193[95]^and_result193[96]^and_result193[97]^and_result193[98]^and_result193[99]^and_result193[100]^and_result193[101]^and_result193[102]^and_result193[103]^and_result193[104]^and_result193[105]^and_result193[106]^and_result193[107]^and_result193[108]^and_result193[109]^and_result193[110]^and_result193[111]^and_result193[112]^and_result193[113]^and_result193[114]^and_result193[115]^and_result193[116]^and_result193[117]^and_result193[118]^and_result193[119]^and_result193[120]^and_result193[121]^and_result193[122]^and_result193[123]^and_result193[124]^and_result193[125]^and_result193[126]^and_result193[127]^and_result193[128]^and_result193[129]^and_result193[130]^and_result193[131]^and_result193[132]^and_result193[133]^and_result193[134]^and_result193[135]^and_result193[136]^and_result193[137]^and_result193[138]^and_result193[139]^and_result193[140]^and_result193[141]^and_result193[142]^and_result193[143]^and_result193[144]^and_result193[145]^and_result193[146]^and_result193[147]^and_result193[148]^and_result193[149]^and_result193[150]^and_result193[151]^and_result193[152]^and_result193[153]^and_result193[154]^and_result193[155]^and_result193[156]^and_result193[157]^and_result193[158]^and_result193[159]^and_result193[160]^and_result193[161]^and_result193[162]^and_result193[163]^and_result193[164]^and_result193[165]^and_result193[166]^and_result193[167]^and_result193[168]^and_result193[169]^and_result193[170]^and_result193[171]^and_result193[172]^and_result193[173]^and_result193[174]^and_result193[175]^and_result193[176]^and_result193[177]^and_result193[178]^and_result193[179]^and_result193[180]^and_result193[181]^and_result193[182]^and_result193[183]^and_result193[184]^and_result193[185]^and_result193[186]^and_result193[187]^and_result193[188]^and_result193[189]^and_result193[190]^and_result193[191]^and_result193[192]^and_result193[193]^and_result193[194]^and_result193[195]^and_result193[196]^and_result193[197]^and_result193[198]^and_result193[199]^and_result193[200]^and_result193[201]^and_result193[202]^and_result193[203]^and_result193[204]^and_result193[205]^and_result193[206]^and_result193[207]^and_result193[208]^and_result193[209]^and_result193[210]^and_result193[211]^and_result193[212]^and_result193[213]^and_result193[214]^and_result193[215]^and_result193[216]^and_result193[217]^and_result193[218]^and_result193[219]^and_result193[220]^and_result193[221]^and_result193[222]^and_result193[223]^and_result193[224]^and_result193[225]^and_result193[226]^and_result193[227]^and_result193[228]^and_result193[229]^and_result193[230]^and_result193[231]^and_result193[232]^and_result193[233]^and_result193[234]^and_result193[235]^and_result193[236]^and_result193[237]^and_result193[238]^and_result193[239]^and_result193[240]^and_result193[241]^and_result193[242]^and_result193[243]^and_result193[244]^and_result193[245]^and_result193[246]^and_result193[247]^and_result193[248]^and_result193[249]^and_result193[250]^and_result193[251]^and_result193[252]^and_result193[253]^and_result193[254];
assign key[194]=and_result194[0]^and_result194[1]^and_result194[2]^and_result194[3]^and_result194[4]^and_result194[5]^and_result194[6]^and_result194[7]^and_result194[8]^and_result194[9]^and_result194[10]^and_result194[11]^and_result194[12]^and_result194[13]^and_result194[14]^and_result194[15]^and_result194[16]^and_result194[17]^and_result194[18]^and_result194[19]^and_result194[20]^and_result194[21]^and_result194[22]^and_result194[23]^and_result194[24]^and_result194[25]^and_result194[26]^and_result194[27]^and_result194[28]^and_result194[29]^and_result194[30]^and_result194[31]^and_result194[32]^and_result194[33]^and_result194[34]^and_result194[35]^and_result194[36]^and_result194[37]^and_result194[38]^and_result194[39]^and_result194[40]^and_result194[41]^and_result194[42]^and_result194[43]^and_result194[44]^and_result194[45]^and_result194[46]^and_result194[47]^and_result194[48]^and_result194[49]^and_result194[50]^and_result194[51]^and_result194[52]^and_result194[53]^and_result194[54]^and_result194[55]^and_result194[56]^and_result194[57]^and_result194[58]^and_result194[59]^and_result194[60]^and_result194[61]^and_result194[62]^and_result194[63]^and_result194[64]^and_result194[65]^and_result194[66]^and_result194[67]^and_result194[68]^and_result194[69]^and_result194[70]^and_result194[71]^and_result194[72]^and_result194[73]^and_result194[74]^and_result194[75]^and_result194[76]^and_result194[77]^and_result194[78]^and_result194[79]^and_result194[80]^and_result194[81]^and_result194[82]^and_result194[83]^and_result194[84]^and_result194[85]^and_result194[86]^and_result194[87]^and_result194[88]^and_result194[89]^and_result194[90]^and_result194[91]^and_result194[92]^and_result194[93]^and_result194[94]^and_result194[95]^and_result194[96]^and_result194[97]^and_result194[98]^and_result194[99]^and_result194[100]^and_result194[101]^and_result194[102]^and_result194[103]^and_result194[104]^and_result194[105]^and_result194[106]^and_result194[107]^and_result194[108]^and_result194[109]^and_result194[110]^and_result194[111]^and_result194[112]^and_result194[113]^and_result194[114]^and_result194[115]^and_result194[116]^and_result194[117]^and_result194[118]^and_result194[119]^and_result194[120]^and_result194[121]^and_result194[122]^and_result194[123]^and_result194[124]^and_result194[125]^and_result194[126]^and_result194[127]^and_result194[128]^and_result194[129]^and_result194[130]^and_result194[131]^and_result194[132]^and_result194[133]^and_result194[134]^and_result194[135]^and_result194[136]^and_result194[137]^and_result194[138]^and_result194[139]^and_result194[140]^and_result194[141]^and_result194[142]^and_result194[143]^and_result194[144]^and_result194[145]^and_result194[146]^and_result194[147]^and_result194[148]^and_result194[149]^and_result194[150]^and_result194[151]^and_result194[152]^and_result194[153]^and_result194[154]^and_result194[155]^and_result194[156]^and_result194[157]^and_result194[158]^and_result194[159]^and_result194[160]^and_result194[161]^and_result194[162]^and_result194[163]^and_result194[164]^and_result194[165]^and_result194[166]^and_result194[167]^and_result194[168]^and_result194[169]^and_result194[170]^and_result194[171]^and_result194[172]^and_result194[173]^and_result194[174]^and_result194[175]^and_result194[176]^and_result194[177]^and_result194[178]^and_result194[179]^and_result194[180]^and_result194[181]^and_result194[182]^and_result194[183]^and_result194[184]^and_result194[185]^and_result194[186]^and_result194[187]^and_result194[188]^and_result194[189]^and_result194[190]^and_result194[191]^and_result194[192]^and_result194[193]^and_result194[194]^and_result194[195]^and_result194[196]^and_result194[197]^and_result194[198]^and_result194[199]^and_result194[200]^and_result194[201]^and_result194[202]^and_result194[203]^and_result194[204]^and_result194[205]^and_result194[206]^and_result194[207]^and_result194[208]^and_result194[209]^and_result194[210]^and_result194[211]^and_result194[212]^and_result194[213]^and_result194[214]^and_result194[215]^and_result194[216]^and_result194[217]^and_result194[218]^and_result194[219]^and_result194[220]^and_result194[221]^and_result194[222]^and_result194[223]^and_result194[224]^and_result194[225]^and_result194[226]^and_result194[227]^and_result194[228]^and_result194[229]^and_result194[230]^and_result194[231]^and_result194[232]^and_result194[233]^and_result194[234]^and_result194[235]^and_result194[236]^and_result194[237]^and_result194[238]^and_result194[239]^and_result194[240]^and_result194[241]^and_result194[242]^and_result194[243]^and_result194[244]^and_result194[245]^and_result194[246]^and_result194[247]^and_result194[248]^and_result194[249]^and_result194[250]^and_result194[251]^and_result194[252]^and_result194[253]^and_result194[254];
assign key[195]=and_result195[0]^and_result195[1]^and_result195[2]^and_result195[3]^and_result195[4]^and_result195[5]^and_result195[6]^and_result195[7]^and_result195[8]^and_result195[9]^and_result195[10]^and_result195[11]^and_result195[12]^and_result195[13]^and_result195[14]^and_result195[15]^and_result195[16]^and_result195[17]^and_result195[18]^and_result195[19]^and_result195[20]^and_result195[21]^and_result195[22]^and_result195[23]^and_result195[24]^and_result195[25]^and_result195[26]^and_result195[27]^and_result195[28]^and_result195[29]^and_result195[30]^and_result195[31]^and_result195[32]^and_result195[33]^and_result195[34]^and_result195[35]^and_result195[36]^and_result195[37]^and_result195[38]^and_result195[39]^and_result195[40]^and_result195[41]^and_result195[42]^and_result195[43]^and_result195[44]^and_result195[45]^and_result195[46]^and_result195[47]^and_result195[48]^and_result195[49]^and_result195[50]^and_result195[51]^and_result195[52]^and_result195[53]^and_result195[54]^and_result195[55]^and_result195[56]^and_result195[57]^and_result195[58]^and_result195[59]^and_result195[60]^and_result195[61]^and_result195[62]^and_result195[63]^and_result195[64]^and_result195[65]^and_result195[66]^and_result195[67]^and_result195[68]^and_result195[69]^and_result195[70]^and_result195[71]^and_result195[72]^and_result195[73]^and_result195[74]^and_result195[75]^and_result195[76]^and_result195[77]^and_result195[78]^and_result195[79]^and_result195[80]^and_result195[81]^and_result195[82]^and_result195[83]^and_result195[84]^and_result195[85]^and_result195[86]^and_result195[87]^and_result195[88]^and_result195[89]^and_result195[90]^and_result195[91]^and_result195[92]^and_result195[93]^and_result195[94]^and_result195[95]^and_result195[96]^and_result195[97]^and_result195[98]^and_result195[99]^and_result195[100]^and_result195[101]^and_result195[102]^and_result195[103]^and_result195[104]^and_result195[105]^and_result195[106]^and_result195[107]^and_result195[108]^and_result195[109]^and_result195[110]^and_result195[111]^and_result195[112]^and_result195[113]^and_result195[114]^and_result195[115]^and_result195[116]^and_result195[117]^and_result195[118]^and_result195[119]^and_result195[120]^and_result195[121]^and_result195[122]^and_result195[123]^and_result195[124]^and_result195[125]^and_result195[126]^and_result195[127]^and_result195[128]^and_result195[129]^and_result195[130]^and_result195[131]^and_result195[132]^and_result195[133]^and_result195[134]^and_result195[135]^and_result195[136]^and_result195[137]^and_result195[138]^and_result195[139]^and_result195[140]^and_result195[141]^and_result195[142]^and_result195[143]^and_result195[144]^and_result195[145]^and_result195[146]^and_result195[147]^and_result195[148]^and_result195[149]^and_result195[150]^and_result195[151]^and_result195[152]^and_result195[153]^and_result195[154]^and_result195[155]^and_result195[156]^and_result195[157]^and_result195[158]^and_result195[159]^and_result195[160]^and_result195[161]^and_result195[162]^and_result195[163]^and_result195[164]^and_result195[165]^and_result195[166]^and_result195[167]^and_result195[168]^and_result195[169]^and_result195[170]^and_result195[171]^and_result195[172]^and_result195[173]^and_result195[174]^and_result195[175]^and_result195[176]^and_result195[177]^and_result195[178]^and_result195[179]^and_result195[180]^and_result195[181]^and_result195[182]^and_result195[183]^and_result195[184]^and_result195[185]^and_result195[186]^and_result195[187]^and_result195[188]^and_result195[189]^and_result195[190]^and_result195[191]^and_result195[192]^and_result195[193]^and_result195[194]^and_result195[195]^and_result195[196]^and_result195[197]^and_result195[198]^and_result195[199]^and_result195[200]^and_result195[201]^and_result195[202]^and_result195[203]^and_result195[204]^and_result195[205]^and_result195[206]^and_result195[207]^and_result195[208]^and_result195[209]^and_result195[210]^and_result195[211]^and_result195[212]^and_result195[213]^and_result195[214]^and_result195[215]^and_result195[216]^and_result195[217]^and_result195[218]^and_result195[219]^and_result195[220]^and_result195[221]^and_result195[222]^and_result195[223]^and_result195[224]^and_result195[225]^and_result195[226]^and_result195[227]^and_result195[228]^and_result195[229]^and_result195[230]^and_result195[231]^and_result195[232]^and_result195[233]^and_result195[234]^and_result195[235]^and_result195[236]^and_result195[237]^and_result195[238]^and_result195[239]^and_result195[240]^and_result195[241]^and_result195[242]^and_result195[243]^and_result195[244]^and_result195[245]^and_result195[246]^and_result195[247]^and_result195[248]^and_result195[249]^and_result195[250]^and_result195[251]^and_result195[252]^and_result195[253]^and_result195[254];
assign key[196]=and_result196[0]^and_result196[1]^and_result196[2]^and_result196[3]^and_result196[4]^and_result196[5]^and_result196[6]^and_result196[7]^and_result196[8]^and_result196[9]^and_result196[10]^and_result196[11]^and_result196[12]^and_result196[13]^and_result196[14]^and_result196[15]^and_result196[16]^and_result196[17]^and_result196[18]^and_result196[19]^and_result196[20]^and_result196[21]^and_result196[22]^and_result196[23]^and_result196[24]^and_result196[25]^and_result196[26]^and_result196[27]^and_result196[28]^and_result196[29]^and_result196[30]^and_result196[31]^and_result196[32]^and_result196[33]^and_result196[34]^and_result196[35]^and_result196[36]^and_result196[37]^and_result196[38]^and_result196[39]^and_result196[40]^and_result196[41]^and_result196[42]^and_result196[43]^and_result196[44]^and_result196[45]^and_result196[46]^and_result196[47]^and_result196[48]^and_result196[49]^and_result196[50]^and_result196[51]^and_result196[52]^and_result196[53]^and_result196[54]^and_result196[55]^and_result196[56]^and_result196[57]^and_result196[58]^and_result196[59]^and_result196[60]^and_result196[61]^and_result196[62]^and_result196[63]^and_result196[64]^and_result196[65]^and_result196[66]^and_result196[67]^and_result196[68]^and_result196[69]^and_result196[70]^and_result196[71]^and_result196[72]^and_result196[73]^and_result196[74]^and_result196[75]^and_result196[76]^and_result196[77]^and_result196[78]^and_result196[79]^and_result196[80]^and_result196[81]^and_result196[82]^and_result196[83]^and_result196[84]^and_result196[85]^and_result196[86]^and_result196[87]^and_result196[88]^and_result196[89]^and_result196[90]^and_result196[91]^and_result196[92]^and_result196[93]^and_result196[94]^and_result196[95]^and_result196[96]^and_result196[97]^and_result196[98]^and_result196[99]^and_result196[100]^and_result196[101]^and_result196[102]^and_result196[103]^and_result196[104]^and_result196[105]^and_result196[106]^and_result196[107]^and_result196[108]^and_result196[109]^and_result196[110]^and_result196[111]^and_result196[112]^and_result196[113]^and_result196[114]^and_result196[115]^and_result196[116]^and_result196[117]^and_result196[118]^and_result196[119]^and_result196[120]^and_result196[121]^and_result196[122]^and_result196[123]^and_result196[124]^and_result196[125]^and_result196[126]^and_result196[127]^and_result196[128]^and_result196[129]^and_result196[130]^and_result196[131]^and_result196[132]^and_result196[133]^and_result196[134]^and_result196[135]^and_result196[136]^and_result196[137]^and_result196[138]^and_result196[139]^and_result196[140]^and_result196[141]^and_result196[142]^and_result196[143]^and_result196[144]^and_result196[145]^and_result196[146]^and_result196[147]^and_result196[148]^and_result196[149]^and_result196[150]^and_result196[151]^and_result196[152]^and_result196[153]^and_result196[154]^and_result196[155]^and_result196[156]^and_result196[157]^and_result196[158]^and_result196[159]^and_result196[160]^and_result196[161]^and_result196[162]^and_result196[163]^and_result196[164]^and_result196[165]^and_result196[166]^and_result196[167]^and_result196[168]^and_result196[169]^and_result196[170]^and_result196[171]^and_result196[172]^and_result196[173]^and_result196[174]^and_result196[175]^and_result196[176]^and_result196[177]^and_result196[178]^and_result196[179]^and_result196[180]^and_result196[181]^and_result196[182]^and_result196[183]^and_result196[184]^and_result196[185]^and_result196[186]^and_result196[187]^and_result196[188]^and_result196[189]^and_result196[190]^and_result196[191]^and_result196[192]^and_result196[193]^and_result196[194]^and_result196[195]^and_result196[196]^and_result196[197]^and_result196[198]^and_result196[199]^and_result196[200]^and_result196[201]^and_result196[202]^and_result196[203]^and_result196[204]^and_result196[205]^and_result196[206]^and_result196[207]^and_result196[208]^and_result196[209]^and_result196[210]^and_result196[211]^and_result196[212]^and_result196[213]^and_result196[214]^and_result196[215]^and_result196[216]^and_result196[217]^and_result196[218]^and_result196[219]^and_result196[220]^and_result196[221]^and_result196[222]^and_result196[223]^and_result196[224]^and_result196[225]^and_result196[226]^and_result196[227]^and_result196[228]^and_result196[229]^and_result196[230]^and_result196[231]^and_result196[232]^and_result196[233]^and_result196[234]^and_result196[235]^and_result196[236]^and_result196[237]^and_result196[238]^and_result196[239]^and_result196[240]^and_result196[241]^and_result196[242]^and_result196[243]^and_result196[244]^and_result196[245]^and_result196[246]^and_result196[247]^and_result196[248]^and_result196[249]^and_result196[250]^and_result196[251]^and_result196[252]^and_result196[253]^and_result196[254];
assign key[197]=and_result197[0]^and_result197[1]^and_result197[2]^and_result197[3]^and_result197[4]^and_result197[5]^and_result197[6]^and_result197[7]^and_result197[8]^and_result197[9]^and_result197[10]^and_result197[11]^and_result197[12]^and_result197[13]^and_result197[14]^and_result197[15]^and_result197[16]^and_result197[17]^and_result197[18]^and_result197[19]^and_result197[20]^and_result197[21]^and_result197[22]^and_result197[23]^and_result197[24]^and_result197[25]^and_result197[26]^and_result197[27]^and_result197[28]^and_result197[29]^and_result197[30]^and_result197[31]^and_result197[32]^and_result197[33]^and_result197[34]^and_result197[35]^and_result197[36]^and_result197[37]^and_result197[38]^and_result197[39]^and_result197[40]^and_result197[41]^and_result197[42]^and_result197[43]^and_result197[44]^and_result197[45]^and_result197[46]^and_result197[47]^and_result197[48]^and_result197[49]^and_result197[50]^and_result197[51]^and_result197[52]^and_result197[53]^and_result197[54]^and_result197[55]^and_result197[56]^and_result197[57]^and_result197[58]^and_result197[59]^and_result197[60]^and_result197[61]^and_result197[62]^and_result197[63]^and_result197[64]^and_result197[65]^and_result197[66]^and_result197[67]^and_result197[68]^and_result197[69]^and_result197[70]^and_result197[71]^and_result197[72]^and_result197[73]^and_result197[74]^and_result197[75]^and_result197[76]^and_result197[77]^and_result197[78]^and_result197[79]^and_result197[80]^and_result197[81]^and_result197[82]^and_result197[83]^and_result197[84]^and_result197[85]^and_result197[86]^and_result197[87]^and_result197[88]^and_result197[89]^and_result197[90]^and_result197[91]^and_result197[92]^and_result197[93]^and_result197[94]^and_result197[95]^and_result197[96]^and_result197[97]^and_result197[98]^and_result197[99]^and_result197[100]^and_result197[101]^and_result197[102]^and_result197[103]^and_result197[104]^and_result197[105]^and_result197[106]^and_result197[107]^and_result197[108]^and_result197[109]^and_result197[110]^and_result197[111]^and_result197[112]^and_result197[113]^and_result197[114]^and_result197[115]^and_result197[116]^and_result197[117]^and_result197[118]^and_result197[119]^and_result197[120]^and_result197[121]^and_result197[122]^and_result197[123]^and_result197[124]^and_result197[125]^and_result197[126]^and_result197[127]^and_result197[128]^and_result197[129]^and_result197[130]^and_result197[131]^and_result197[132]^and_result197[133]^and_result197[134]^and_result197[135]^and_result197[136]^and_result197[137]^and_result197[138]^and_result197[139]^and_result197[140]^and_result197[141]^and_result197[142]^and_result197[143]^and_result197[144]^and_result197[145]^and_result197[146]^and_result197[147]^and_result197[148]^and_result197[149]^and_result197[150]^and_result197[151]^and_result197[152]^and_result197[153]^and_result197[154]^and_result197[155]^and_result197[156]^and_result197[157]^and_result197[158]^and_result197[159]^and_result197[160]^and_result197[161]^and_result197[162]^and_result197[163]^and_result197[164]^and_result197[165]^and_result197[166]^and_result197[167]^and_result197[168]^and_result197[169]^and_result197[170]^and_result197[171]^and_result197[172]^and_result197[173]^and_result197[174]^and_result197[175]^and_result197[176]^and_result197[177]^and_result197[178]^and_result197[179]^and_result197[180]^and_result197[181]^and_result197[182]^and_result197[183]^and_result197[184]^and_result197[185]^and_result197[186]^and_result197[187]^and_result197[188]^and_result197[189]^and_result197[190]^and_result197[191]^and_result197[192]^and_result197[193]^and_result197[194]^and_result197[195]^and_result197[196]^and_result197[197]^and_result197[198]^and_result197[199]^and_result197[200]^and_result197[201]^and_result197[202]^and_result197[203]^and_result197[204]^and_result197[205]^and_result197[206]^and_result197[207]^and_result197[208]^and_result197[209]^and_result197[210]^and_result197[211]^and_result197[212]^and_result197[213]^and_result197[214]^and_result197[215]^and_result197[216]^and_result197[217]^and_result197[218]^and_result197[219]^and_result197[220]^and_result197[221]^and_result197[222]^and_result197[223]^and_result197[224]^and_result197[225]^and_result197[226]^and_result197[227]^and_result197[228]^and_result197[229]^and_result197[230]^and_result197[231]^and_result197[232]^and_result197[233]^and_result197[234]^and_result197[235]^and_result197[236]^and_result197[237]^and_result197[238]^and_result197[239]^and_result197[240]^and_result197[241]^and_result197[242]^and_result197[243]^and_result197[244]^and_result197[245]^and_result197[246]^and_result197[247]^and_result197[248]^and_result197[249]^and_result197[250]^and_result197[251]^and_result197[252]^and_result197[253]^and_result197[254];
assign key[198]=and_result198[0]^and_result198[1]^and_result198[2]^and_result198[3]^and_result198[4]^and_result198[5]^and_result198[6]^and_result198[7]^and_result198[8]^and_result198[9]^and_result198[10]^and_result198[11]^and_result198[12]^and_result198[13]^and_result198[14]^and_result198[15]^and_result198[16]^and_result198[17]^and_result198[18]^and_result198[19]^and_result198[20]^and_result198[21]^and_result198[22]^and_result198[23]^and_result198[24]^and_result198[25]^and_result198[26]^and_result198[27]^and_result198[28]^and_result198[29]^and_result198[30]^and_result198[31]^and_result198[32]^and_result198[33]^and_result198[34]^and_result198[35]^and_result198[36]^and_result198[37]^and_result198[38]^and_result198[39]^and_result198[40]^and_result198[41]^and_result198[42]^and_result198[43]^and_result198[44]^and_result198[45]^and_result198[46]^and_result198[47]^and_result198[48]^and_result198[49]^and_result198[50]^and_result198[51]^and_result198[52]^and_result198[53]^and_result198[54]^and_result198[55]^and_result198[56]^and_result198[57]^and_result198[58]^and_result198[59]^and_result198[60]^and_result198[61]^and_result198[62]^and_result198[63]^and_result198[64]^and_result198[65]^and_result198[66]^and_result198[67]^and_result198[68]^and_result198[69]^and_result198[70]^and_result198[71]^and_result198[72]^and_result198[73]^and_result198[74]^and_result198[75]^and_result198[76]^and_result198[77]^and_result198[78]^and_result198[79]^and_result198[80]^and_result198[81]^and_result198[82]^and_result198[83]^and_result198[84]^and_result198[85]^and_result198[86]^and_result198[87]^and_result198[88]^and_result198[89]^and_result198[90]^and_result198[91]^and_result198[92]^and_result198[93]^and_result198[94]^and_result198[95]^and_result198[96]^and_result198[97]^and_result198[98]^and_result198[99]^and_result198[100]^and_result198[101]^and_result198[102]^and_result198[103]^and_result198[104]^and_result198[105]^and_result198[106]^and_result198[107]^and_result198[108]^and_result198[109]^and_result198[110]^and_result198[111]^and_result198[112]^and_result198[113]^and_result198[114]^and_result198[115]^and_result198[116]^and_result198[117]^and_result198[118]^and_result198[119]^and_result198[120]^and_result198[121]^and_result198[122]^and_result198[123]^and_result198[124]^and_result198[125]^and_result198[126]^and_result198[127]^and_result198[128]^and_result198[129]^and_result198[130]^and_result198[131]^and_result198[132]^and_result198[133]^and_result198[134]^and_result198[135]^and_result198[136]^and_result198[137]^and_result198[138]^and_result198[139]^and_result198[140]^and_result198[141]^and_result198[142]^and_result198[143]^and_result198[144]^and_result198[145]^and_result198[146]^and_result198[147]^and_result198[148]^and_result198[149]^and_result198[150]^and_result198[151]^and_result198[152]^and_result198[153]^and_result198[154]^and_result198[155]^and_result198[156]^and_result198[157]^and_result198[158]^and_result198[159]^and_result198[160]^and_result198[161]^and_result198[162]^and_result198[163]^and_result198[164]^and_result198[165]^and_result198[166]^and_result198[167]^and_result198[168]^and_result198[169]^and_result198[170]^and_result198[171]^and_result198[172]^and_result198[173]^and_result198[174]^and_result198[175]^and_result198[176]^and_result198[177]^and_result198[178]^and_result198[179]^and_result198[180]^and_result198[181]^and_result198[182]^and_result198[183]^and_result198[184]^and_result198[185]^and_result198[186]^and_result198[187]^and_result198[188]^and_result198[189]^and_result198[190]^and_result198[191]^and_result198[192]^and_result198[193]^and_result198[194]^and_result198[195]^and_result198[196]^and_result198[197]^and_result198[198]^and_result198[199]^and_result198[200]^and_result198[201]^and_result198[202]^and_result198[203]^and_result198[204]^and_result198[205]^and_result198[206]^and_result198[207]^and_result198[208]^and_result198[209]^and_result198[210]^and_result198[211]^and_result198[212]^and_result198[213]^and_result198[214]^and_result198[215]^and_result198[216]^and_result198[217]^and_result198[218]^and_result198[219]^and_result198[220]^and_result198[221]^and_result198[222]^and_result198[223]^and_result198[224]^and_result198[225]^and_result198[226]^and_result198[227]^and_result198[228]^and_result198[229]^and_result198[230]^and_result198[231]^and_result198[232]^and_result198[233]^and_result198[234]^and_result198[235]^and_result198[236]^and_result198[237]^and_result198[238]^and_result198[239]^and_result198[240]^and_result198[241]^and_result198[242]^and_result198[243]^and_result198[244]^and_result198[245]^and_result198[246]^and_result198[247]^and_result198[248]^and_result198[249]^and_result198[250]^and_result198[251]^and_result198[252]^and_result198[253]^and_result198[254];
assign key[199]=and_result199[0]^and_result199[1]^and_result199[2]^and_result199[3]^and_result199[4]^and_result199[5]^and_result199[6]^and_result199[7]^and_result199[8]^and_result199[9]^and_result199[10]^and_result199[11]^and_result199[12]^and_result199[13]^and_result199[14]^and_result199[15]^and_result199[16]^and_result199[17]^and_result199[18]^and_result199[19]^and_result199[20]^and_result199[21]^and_result199[22]^and_result199[23]^and_result199[24]^and_result199[25]^and_result199[26]^and_result199[27]^and_result199[28]^and_result199[29]^and_result199[30]^and_result199[31]^and_result199[32]^and_result199[33]^and_result199[34]^and_result199[35]^and_result199[36]^and_result199[37]^and_result199[38]^and_result199[39]^and_result199[40]^and_result199[41]^and_result199[42]^and_result199[43]^and_result199[44]^and_result199[45]^and_result199[46]^and_result199[47]^and_result199[48]^and_result199[49]^and_result199[50]^and_result199[51]^and_result199[52]^and_result199[53]^and_result199[54]^and_result199[55]^and_result199[56]^and_result199[57]^and_result199[58]^and_result199[59]^and_result199[60]^and_result199[61]^and_result199[62]^and_result199[63]^and_result199[64]^and_result199[65]^and_result199[66]^and_result199[67]^and_result199[68]^and_result199[69]^and_result199[70]^and_result199[71]^and_result199[72]^and_result199[73]^and_result199[74]^and_result199[75]^and_result199[76]^and_result199[77]^and_result199[78]^and_result199[79]^and_result199[80]^and_result199[81]^and_result199[82]^and_result199[83]^and_result199[84]^and_result199[85]^and_result199[86]^and_result199[87]^and_result199[88]^and_result199[89]^and_result199[90]^and_result199[91]^and_result199[92]^and_result199[93]^and_result199[94]^and_result199[95]^and_result199[96]^and_result199[97]^and_result199[98]^and_result199[99]^and_result199[100]^and_result199[101]^and_result199[102]^and_result199[103]^and_result199[104]^and_result199[105]^and_result199[106]^and_result199[107]^and_result199[108]^and_result199[109]^and_result199[110]^and_result199[111]^and_result199[112]^and_result199[113]^and_result199[114]^and_result199[115]^and_result199[116]^and_result199[117]^and_result199[118]^and_result199[119]^and_result199[120]^and_result199[121]^and_result199[122]^and_result199[123]^and_result199[124]^and_result199[125]^and_result199[126]^and_result199[127]^and_result199[128]^and_result199[129]^and_result199[130]^and_result199[131]^and_result199[132]^and_result199[133]^and_result199[134]^and_result199[135]^and_result199[136]^and_result199[137]^and_result199[138]^and_result199[139]^and_result199[140]^and_result199[141]^and_result199[142]^and_result199[143]^and_result199[144]^and_result199[145]^and_result199[146]^and_result199[147]^and_result199[148]^and_result199[149]^and_result199[150]^and_result199[151]^and_result199[152]^and_result199[153]^and_result199[154]^and_result199[155]^and_result199[156]^and_result199[157]^and_result199[158]^and_result199[159]^and_result199[160]^and_result199[161]^and_result199[162]^and_result199[163]^and_result199[164]^and_result199[165]^and_result199[166]^and_result199[167]^and_result199[168]^and_result199[169]^and_result199[170]^and_result199[171]^and_result199[172]^and_result199[173]^and_result199[174]^and_result199[175]^and_result199[176]^and_result199[177]^and_result199[178]^and_result199[179]^and_result199[180]^and_result199[181]^and_result199[182]^and_result199[183]^and_result199[184]^and_result199[185]^and_result199[186]^and_result199[187]^and_result199[188]^and_result199[189]^and_result199[190]^and_result199[191]^and_result199[192]^and_result199[193]^and_result199[194]^and_result199[195]^and_result199[196]^and_result199[197]^and_result199[198]^and_result199[199]^and_result199[200]^and_result199[201]^and_result199[202]^and_result199[203]^and_result199[204]^and_result199[205]^and_result199[206]^and_result199[207]^and_result199[208]^and_result199[209]^and_result199[210]^and_result199[211]^and_result199[212]^and_result199[213]^and_result199[214]^and_result199[215]^and_result199[216]^and_result199[217]^and_result199[218]^and_result199[219]^and_result199[220]^and_result199[221]^and_result199[222]^and_result199[223]^and_result199[224]^and_result199[225]^and_result199[226]^and_result199[227]^and_result199[228]^and_result199[229]^and_result199[230]^and_result199[231]^and_result199[232]^and_result199[233]^and_result199[234]^and_result199[235]^and_result199[236]^and_result199[237]^and_result199[238]^and_result199[239]^and_result199[240]^and_result199[241]^and_result199[242]^and_result199[243]^and_result199[244]^and_result199[245]^and_result199[246]^and_result199[247]^and_result199[248]^and_result199[249]^and_result199[250]^and_result199[251]^and_result199[252]^and_result199[253]^and_result199[254];
assign key[200]=and_result200[0]^and_result200[1]^and_result200[2]^and_result200[3]^and_result200[4]^and_result200[5]^and_result200[6]^and_result200[7]^and_result200[8]^and_result200[9]^and_result200[10]^and_result200[11]^and_result200[12]^and_result200[13]^and_result200[14]^and_result200[15]^and_result200[16]^and_result200[17]^and_result200[18]^and_result200[19]^and_result200[20]^and_result200[21]^and_result200[22]^and_result200[23]^and_result200[24]^and_result200[25]^and_result200[26]^and_result200[27]^and_result200[28]^and_result200[29]^and_result200[30]^and_result200[31]^and_result200[32]^and_result200[33]^and_result200[34]^and_result200[35]^and_result200[36]^and_result200[37]^and_result200[38]^and_result200[39]^and_result200[40]^and_result200[41]^and_result200[42]^and_result200[43]^and_result200[44]^and_result200[45]^and_result200[46]^and_result200[47]^and_result200[48]^and_result200[49]^and_result200[50]^and_result200[51]^and_result200[52]^and_result200[53]^and_result200[54]^and_result200[55]^and_result200[56]^and_result200[57]^and_result200[58]^and_result200[59]^and_result200[60]^and_result200[61]^and_result200[62]^and_result200[63]^and_result200[64]^and_result200[65]^and_result200[66]^and_result200[67]^and_result200[68]^and_result200[69]^and_result200[70]^and_result200[71]^and_result200[72]^and_result200[73]^and_result200[74]^and_result200[75]^and_result200[76]^and_result200[77]^and_result200[78]^and_result200[79]^and_result200[80]^and_result200[81]^and_result200[82]^and_result200[83]^and_result200[84]^and_result200[85]^and_result200[86]^and_result200[87]^and_result200[88]^and_result200[89]^and_result200[90]^and_result200[91]^and_result200[92]^and_result200[93]^and_result200[94]^and_result200[95]^and_result200[96]^and_result200[97]^and_result200[98]^and_result200[99]^and_result200[100]^and_result200[101]^and_result200[102]^and_result200[103]^and_result200[104]^and_result200[105]^and_result200[106]^and_result200[107]^and_result200[108]^and_result200[109]^and_result200[110]^and_result200[111]^and_result200[112]^and_result200[113]^and_result200[114]^and_result200[115]^and_result200[116]^and_result200[117]^and_result200[118]^and_result200[119]^and_result200[120]^and_result200[121]^and_result200[122]^and_result200[123]^and_result200[124]^and_result200[125]^and_result200[126]^and_result200[127]^and_result200[128]^and_result200[129]^and_result200[130]^and_result200[131]^and_result200[132]^and_result200[133]^and_result200[134]^and_result200[135]^and_result200[136]^and_result200[137]^and_result200[138]^and_result200[139]^and_result200[140]^and_result200[141]^and_result200[142]^and_result200[143]^and_result200[144]^and_result200[145]^and_result200[146]^and_result200[147]^and_result200[148]^and_result200[149]^and_result200[150]^and_result200[151]^and_result200[152]^and_result200[153]^and_result200[154]^and_result200[155]^and_result200[156]^and_result200[157]^and_result200[158]^and_result200[159]^and_result200[160]^and_result200[161]^and_result200[162]^and_result200[163]^and_result200[164]^and_result200[165]^and_result200[166]^and_result200[167]^and_result200[168]^and_result200[169]^and_result200[170]^and_result200[171]^and_result200[172]^and_result200[173]^and_result200[174]^and_result200[175]^and_result200[176]^and_result200[177]^and_result200[178]^and_result200[179]^and_result200[180]^and_result200[181]^and_result200[182]^and_result200[183]^and_result200[184]^and_result200[185]^and_result200[186]^and_result200[187]^and_result200[188]^and_result200[189]^and_result200[190]^and_result200[191]^and_result200[192]^and_result200[193]^and_result200[194]^and_result200[195]^and_result200[196]^and_result200[197]^and_result200[198]^and_result200[199]^and_result200[200]^and_result200[201]^and_result200[202]^and_result200[203]^and_result200[204]^and_result200[205]^and_result200[206]^and_result200[207]^and_result200[208]^and_result200[209]^and_result200[210]^and_result200[211]^and_result200[212]^and_result200[213]^and_result200[214]^and_result200[215]^and_result200[216]^and_result200[217]^and_result200[218]^and_result200[219]^and_result200[220]^and_result200[221]^and_result200[222]^and_result200[223]^and_result200[224]^and_result200[225]^and_result200[226]^and_result200[227]^and_result200[228]^and_result200[229]^and_result200[230]^and_result200[231]^and_result200[232]^and_result200[233]^and_result200[234]^and_result200[235]^and_result200[236]^and_result200[237]^and_result200[238]^and_result200[239]^and_result200[240]^and_result200[241]^and_result200[242]^and_result200[243]^and_result200[244]^and_result200[245]^and_result200[246]^and_result200[247]^and_result200[248]^and_result200[249]^and_result200[250]^and_result200[251]^and_result200[252]^and_result200[253]^and_result200[254];
assign key[201]=and_result201[0]^and_result201[1]^and_result201[2]^and_result201[3]^and_result201[4]^and_result201[5]^and_result201[6]^and_result201[7]^and_result201[8]^and_result201[9]^and_result201[10]^and_result201[11]^and_result201[12]^and_result201[13]^and_result201[14]^and_result201[15]^and_result201[16]^and_result201[17]^and_result201[18]^and_result201[19]^and_result201[20]^and_result201[21]^and_result201[22]^and_result201[23]^and_result201[24]^and_result201[25]^and_result201[26]^and_result201[27]^and_result201[28]^and_result201[29]^and_result201[30]^and_result201[31]^and_result201[32]^and_result201[33]^and_result201[34]^and_result201[35]^and_result201[36]^and_result201[37]^and_result201[38]^and_result201[39]^and_result201[40]^and_result201[41]^and_result201[42]^and_result201[43]^and_result201[44]^and_result201[45]^and_result201[46]^and_result201[47]^and_result201[48]^and_result201[49]^and_result201[50]^and_result201[51]^and_result201[52]^and_result201[53]^and_result201[54]^and_result201[55]^and_result201[56]^and_result201[57]^and_result201[58]^and_result201[59]^and_result201[60]^and_result201[61]^and_result201[62]^and_result201[63]^and_result201[64]^and_result201[65]^and_result201[66]^and_result201[67]^and_result201[68]^and_result201[69]^and_result201[70]^and_result201[71]^and_result201[72]^and_result201[73]^and_result201[74]^and_result201[75]^and_result201[76]^and_result201[77]^and_result201[78]^and_result201[79]^and_result201[80]^and_result201[81]^and_result201[82]^and_result201[83]^and_result201[84]^and_result201[85]^and_result201[86]^and_result201[87]^and_result201[88]^and_result201[89]^and_result201[90]^and_result201[91]^and_result201[92]^and_result201[93]^and_result201[94]^and_result201[95]^and_result201[96]^and_result201[97]^and_result201[98]^and_result201[99]^and_result201[100]^and_result201[101]^and_result201[102]^and_result201[103]^and_result201[104]^and_result201[105]^and_result201[106]^and_result201[107]^and_result201[108]^and_result201[109]^and_result201[110]^and_result201[111]^and_result201[112]^and_result201[113]^and_result201[114]^and_result201[115]^and_result201[116]^and_result201[117]^and_result201[118]^and_result201[119]^and_result201[120]^and_result201[121]^and_result201[122]^and_result201[123]^and_result201[124]^and_result201[125]^and_result201[126]^and_result201[127]^and_result201[128]^and_result201[129]^and_result201[130]^and_result201[131]^and_result201[132]^and_result201[133]^and_result201[134]^and_result201[135]^and_result201[136]^and_result201[137]^and_result201[138]^and_result201[139]^and_result201[140]^and_result201[141]^and_result201[142]^and_result201[143]^and_result201[144]^and_result201[145]^and_result201[146]^and_result201[147]^and_result201[148]^and_result201[149]^and_result201[150]^and_result201[151]^and_result201[152]^and_result201[153]^and_result201[154]^and_result201[155]^and_result201[156]^and_result201[157]^and_result201[158]^and_result201[159]^and_result201[160]^and_result201[161]^and_result201[162]^and_result201[163]^and_result201[164]^and_result201[165]^and_result201[166]^and_result201[167]^and_result201[168]^and_result201[169]^and_result201[170]^and_result201[171]^and_result201[172]^and_result201[173]^and_result201[174]^and_result201[175]^and_result201[176]^and_result201[177]^and_result201[178]^and_result201[179]^and_result201[180]^and_result201[181]^and_result201[182]^and_result201[183]^and_result201[184]^and_result201[185]^and_result201[186]^and_result201[187]^and_result201[188]^and_result201[189]^and_result201[190]^and_result201[191]^and_result201[192]^and_result201[193]^and_result201[194]^and_result201[195]^and_result201[196]^and_result201[197]^and_result201[198]^and_result201[199]^and_result201[200]^and_result201[201]^and_result201[202]^and_result201[203]^and_result201[204]^and_result201[205]^and_result201[206]^and_result201[207]^and_result201[208]^and_result201[209]^and_result201[210]^and_result201[211]^and_result201[212]^and_result201[213]^and_result201[214]^and_result201[215]^and_result201[216]^and_result201[217]^and_result201[218]^and_result201[219]^and_result201[220]^and_result201[221]^and_result201[222]^and_result201[223]^and_result201[224]^and_result201[225]^and_result201[226]^and_result201[227]^and_result201[228]^and_result201[229]^and_result201[230]^and_result201[231]^and_result201[232]^and_result201[233]^and_result201[234]^and_result201[235]^and_result201[236]^and_result201[237]^and_result201[238]^and_result201[239]^and_result201[240]^and_result201[241]^and_result201[242]^and_result201[243]^and_result201[244]^and_result201[245]^and_result201[246]^and_result201[247]^and_result201[248]^and_result201[249]^and_result201[250]^and_result201[251]^and_result201[252]^and_result201[253]^and_result201[254];
assign key[202]=and_result202[0]^and_result202[1]^and_result202[2]^and_result202[3]^and_result202[4]^and_result202[5]^and_result202[6]^and_result202[7]^and_result202[8]^and_result202[9]^and_result202[10]^and_result202[11]^and_result202[12]^and_result202[13]^and_result202[14]^and_result202[15]^and_result202[16]^and_result202[17]^and_result202[18]^and_result202[19]^and_result202[20]^and_result202[21]^and_result202[22]^and_result202[23]^and_result202[24]^and_result202[25]^and_result202[26]^and_result202[27]^and_result202[28]^and_result202[29]^and_result202[30]^and_result202[31]^and_result202[32]^and_result202[33]^and_result202[34]^and_result202[35]^and_result202[36]^and_result202[37]^and_result202[38]^and_result202[39]^and_result202[40]^and_result202[41]^and_result202[42]^and_result202[43]^and_result202[44]^and_result202[45]^and_result202[46]^and_result202[47]^and_result202[48]^and_result202[49]^and_result202[50]^and_result202[51]^and_result202[52]^and_result202[53]^and_result202[54]^and_result202[55]^and_result202[56]^and_result202[57]^and_result202[58]^and_result202[59]^and_result202[60]^and_result202[61]^and_result202[62]^and_result202[63]^and_result202[64]^and_result202[65]^and_result202[66]^and_result202[67]^and_result202[68]^and_result202[69]^and_result202[70]^and_result202[71]^and_result202[72]^and_result202[73]^and_result202[74]^and_result202[75]^and_result202[76]^and_result202[77]^and_result202[78]^and_result202[79]^and_result202[80]^and_result202[81]^and_result202[82]^and_result202[83]^and_result202[84]^and_result202[85]^and_result202[86]^and_result202[87]^and_result202[88]^and_result202[89]^and_result202[90]^and_result202[91]^and_result202[92]^and_result202[93]^and_result202[94]^and_result202[95]^and_result202[96]^and_result202[97]^and_result202[98]^and_result202[99]^and_result202[100]^and_result202[101]^and_result202[102]^and_result202[103]^and_result202[104]^and_result202[105]^and_result202[106]^and_result202[107]^and_result202[108]^and_result202[109]^and_result202[110]^and_result202[111]^and_result202[112]^and_result202[113]^and_result202[114]^and_result202[115]^and_result202[116]^and_result202[117]^and_result202[118]^and_result202[119]^and_result202[120]^and_result202[121]^and_result202[122]^and_result202[123]^and_result202[124]^and_result202[125]^and_result202[126]^and_result202[127]^and_result202[128]^and_result202[129]^and_result202[130]^and_result202[131]^and_result202[132]^and_result202[133]^and_result202[134]^and_result202[135]^and_result202[136]^and_result202[137]^and_result202[138]^and_result202[139]^and_result202[140]^and_result202[141]^and_result202[142]^and_result202[143]^and_result202[144]^and_result202[145]^and_result202[146]^and_result202[147]^and_result202[148]^and_result202[149]^and_result202[150]^and_result202[151]^and_result202[152]^and_result202[153]^and_result202[154]^and_result202[155]^and_result202[156]^and_result202[157]^and_result202[158]^and_result202[159]^and_result202[160]^and_result202[161]^and_result202[162]^and_result202[163]^and_result202[164]^and_result202[165]^and_result202[166]^and_result202[167]^and_result202[168]^and_result202[169]^and_result202[170]^and_result202[171]^and_result202[172]^and_result202[173]^and_result202[174]^and_result202[175]^and_result202[176]^and_result202[177]^and_result202[178]^and_result202[179]^and_result202[180]^and_result202[181]^and_result202[182]^and_result202[183]^and_result202[184]^and_result202[185]^and_result202[186]^and_result202[187]^and_result202[188]^and_result202[189]^and_result202[190]^and_result202[191]^and_result202[192]^and_result202[193]^and_result202[194]^and_result202[195]^and_result202[196]^and_result202[197]^and_result202[198]^and_result202[199]^and_result202[200]^and_result202[201]^and_result202[202]^and_result202[203]^and_result202[204]^and_result202[205]^and_result202[206]^and_result202[207]^and_result202[208]^and_result202[209]^and_result202[210]^and_result202[211]^and_result202[212]^and_result202[213]^and_result202[214]^and_result202[215]^and_result202[216]^and_result202[217]^and_result202[218]^and_result202[219]^and_result202[220]^and_result202[221]^and_result202[222]^and_result202[223]^and_result202[224]^and_result202[225]^and_result202[226]^and_result202[227]^and_result202[228]^and_result202[229]^and_result202[230]^and_result202[231]^and_result202[232]^and_result202[233]^and_result202[234]^and_result202[235]^and_result202[236]^and_result202[237]^and_result202[238]^and_result202[239]^and_result202[240]^and_result202[241]^and_result202[242]^and_result202[243]^and_result202[244]^and_result202[245]^and_result202[246]^and_result202[247]^and_result202[248]^and_result202[249]^and_result202[250]^and_result202[251]^and_result202[252]^and_result202[253]^and_result202[254];
assign key[203]=and_result203[0]^and_result203[1]^and_result203[2]^and_result203[3]^and_result203[4]^and_result203[5]^and_result203[6]^and_result203[7]^and_result203[8]^and_result203[9]^and_result203[10]^and_result203[11]^and_result203[12]^and_result203[13]^and_result203[14]^and_result203[15]^and_result203[16]^and_result203[17]^and_result203[18]^and_result203[19]^and_result203[20]^and_result203[21]^and_result203[22]^and_result203[23]^and_result203[24]^and_result203[25]^and_result203[26]^and_result203[27]^and_result203[28]^and_result203[29]^and_result203[30]^and_result203[31]^and_result203[32]^and_result203[33]^and_result203[34]^and_result203[35]^and_result203[36]^and_result203[37]^and_result203[38]^and_result203[39]^and_result203[40]^and_result203[41]^and_result203[42]^and_result203[43]^and_result203[44]^and_result203[45]^and_result203[46]^and_result203[47]^and_result203[48]^and_result203[49]^and_result203[50]^and_result203[51]^and_result203[52]^and_result203[53]^and_result203[54]^and_result203[55]^and_result203[56]^and_result203[57]^and_result203[58]^and_result203[59]^and_result203[60]^and_result203[61]^and_result203[62]^and_result203[63]^and_result203[64]^and_result203[65]^and_result203[66]^and_result203[67]^and_result203[68]^and_result203[69]^and_result203[70]^and_result203[71]^and_result203[72]^and_result203[73]^and_result203[74]^and_result203[75]^and_result203[76]^and_result203[77]^and_result203[78]^and_result203[79]^and_result203[80]^and_result203[81]^and_result203[82]^and_result203[83]^and_result203[84]^and_result203[85]^and_result203[86]^and_result203[87]^and_result203[88]^and_result203[89]^and_result203[90]^and_result203[91]^and_result203[92]^and_result203[93]^and_result203[94]^and_result203[95]^and_result203[96]^and_result203[97]^and_result203[98]^and_result203[99]^and_result203[100]^and_result203[101]^and_result203[102]^and_result203[103]^and_result203[104]^and_result203[105]^and_result203[106]^and_result203[107]^and_result203[108]^and_result203[109]^and_result203[110]^and_result203[111]^and_result203[112]^and_result203[113]^and_result203[114]^and_result203[115]^and_result203[116]^and_result203[117]^and_result203[118]^and_result203[119]^and_result203[120]^and_result203[121]^and_result203[122]^and_result203[123]^and_result203[124]^and_result203[125]^and_result203[126]^and_result203[127]^and_result203[128]^and_result203[129]^and_result203[130]^and_result203[131]^and_result203[132]^and_result203[133]^and_result203[134]^and_result203[135]^and_result203[136]^and_result203[137]^and_result203[138]^and_result203[139]^and_result203[140]^and_result203[141]^and_result203[142]^and_result203[143]^and_result203[144]^and_result203[145]^and_result203[146]^and_result203[147]^and_result203[148]^and_result203[149]^and_result203[150]^and_result203[151]^and_result203[152]^and_result203[153]^and_result203[154]^and_result203[155]^and_result203[156]^and_result203[157]^and_result203[158]^and_result203[159]^and_result203[160]^and_result203[161]^and_result203[162]^and_result203[163]^and_result203[164]^and_result203[165]^and_result203[166]^and_result203[167]^and_result203[168]^and_result203[169]^and_result203[170]^and_result203[171]^and_result203[172]^and_result203[173]^and_result203[174]^and_result203[175]^and_result203[176]^and_result203[177]^and_result203[178]^and_result203[179]^and_result203[180]^and_result203[181]^and_result203[182]^and_result203[183]^and_result203[184]^and_result203[185]^and_result203[186]^and_result203[187]^and_result203[188]^and_result203[189]^and_result203[190]^and_result203[191]^and_result203[192]^and_result203[193]^and_result203[194]^and_result203[195]^and_result203[196]^and_result203[197]^and_result203[198]^and_result203[199]^and_result203[200]^and_result203[201]^and_result203[202]^and_result203[203]^and_result203[204]^and_result203[205]^and_result203[206]^and_result203[207]^and_result203[208]^and_result203[209]^and_result203[210]^and_result203[211]^and_result203[212]^and_result203[213]^and_result203[214]^and_result203[215]^and_result203[216]^and_result203[217]^and_result203[218]^and_result203[219]^and_result203[220]^and_result203[221]^and_result203[222]^and_result203[223]^and_result203[224]^and_result203[225]^and_result203[226]^and_result203[227]^and_result203[228]^and_result203[229]^and_result203[230]^and_result203[231]^and_result203[232]^and_result203[233]^and_result203[234]^and_result203[235]^and_result203[236]^and_result203[237]^and_result203[238]^and_result203[239]^and_result203[240]^and_result203[241]^and_result203[242]^and_result203[243]^and_result203[244]^and_result203[245]^and_result203[246]^and_result203[247]^and_result203[248]^and_result203[249]^and_result203[250]^and_result203[251]^and_result203[252]^and_result203[253]^and_result203[254];
assign key[204]=and_result204[0]^and_result204[1]^and_result204[2]^and_result204[3]^and_result204[4]^and_result204[5]^and_result204[6]^and_result204[7]^and_result204[8]^and_result204[9]^and_result204[10]^and_result204[11]^and_result204[12]^and_result204[13]^and_result204[14]^and_result204[15]^and_result204[16]^and_result204[17]^and_result204[18]^and_result204[19]^and_result204[20]^and_result204[21]^and_result204[22]^and_result204[23]^and_result204[24]^and_result204[25]^and_result204[26]^and_result204[27]^and_result204[28]^and_result204[29]^and_result204[30]^and_result204[31]^and_result204[32]^and_result204[33]^and_result204[34]^and_result204[35]^and_result204[36]^and_result204[37]^and_result204[38]^and_result204[39]^and_result204[40]^and_result204[41]^and_result204[42]^and_result204[43]^and_result204[44]^and_result204[45]^and_result204[46]^and_result204[47]^and_result204[48]^and_result204[49]^and_result204[50]^and_result204[51]^and_result204[52]^and_result204[53]^and_result204[54]^and_result204[55]^and_result204[56]^and_result204[57]^and_result204[58]^and_result204[59]^and_result204[60]^and_result204[61]^and_result204[62]^and_result204[63]^and_result204[64]^and_result204[65]^and_result204[66]^and_result204[67]^and_result204[68]^and_result204[69]^and_result204[70]^and_result204[71]^and_result204[72]^and_result204[73]^and_result204[74]^and_result204[75]^and_result204[76]^and_result204[77]^and_result204[78]^and_result204[79]^and_result204[80]^and_result204[81]^and_result204[82]^and_result204[83]^and_result204[84]^and_result204[85]^and_result204[86]^and_result204[87]^and_result204[88]^and_result204[89]^and_result204[90]^and_result204[91]^and_result204[92]^and_result204[93]^and_result204[94]^and_result204[95]^and_result204[96]^and_result204[97]^and_result204[98]^and_result204[99]^and_result204[100]^and_result204[101]^and_result204[102]^and_result204[103]^and_result204[104]^and_result204[105]^and_result204[106]^and_result204[107]^and_result204[108]^and_result204[109]^and_result204[110]^and_result204[111]^and_result204[112]^and_result204[113]^and_result204[114]^and_result204[115]^and_result204[116]^and_result204[117]^and_result204[118]^and_result204[119]^and_result204[120]^and_result204[121]^and_result204[122]^and_result204[123]^and_result204[124]^and_result204[125]^and_result204[126]^and_result204[127]^and_result204[128]^and_result204[129]^and_result204[130]^and_result204[131]^and_result204[132]^and_result204[133]^and_result204[134]^and_result204[135]^and_result204[136]^and_result204[137]^and_result204[138]^and_result204[139]^and_result204[140]^and_result204[141]^and_result204[142]^and_result204[143]^and_result204[144]^and_result204[145]^and_result204[146]^and_result204[147]^and_result204[148]^and_result204[149]^and_result204[150]^and_result204[151]^and_result204[152]^and_result204[153]^and_result204[154]^and_result204[155]^and_result204[156]^and_result204[157]^and_result204[158]^and_result204[159]^and_result204[160]^and_result204[161]^and_result204[162]^and_result204[163]^and_result204[164]^and_result204[165]^and_result204[166]^and_result204[167]^and_result204[168]^and_result204[169]^and_result204[170]^and_result204[171]^and_result204[172]^and_result204[173]^and_result204[174]^and_result204[175]^and_result204[176]^and_result204[177]^and_result204[178]^and_result204[179]^and_result204[180]^and_result204[181]^and_result204[182]^and_result204[183]^and_result204[184]^and_result204[185]^and_result204[186]^and_result204[187]^and_result204[188]^and_result204[189]^and_result204[190]^and_result204[191]^and_result204[192]^and_result204[193]^and_result204[194]^and_result204[195]^and_result204[196]^and_result204[197]^and_result204[198]^and_result204[199]^and_result204[200]^and_result204[201]^and_result204[202]^and_result204[203]^and_result204[204]^and_result204[205]^and_result204[206]^and_result204[207]^and_result204[208]^and_result204[209]^and_result204[210]^and_result204[211]^and_result204[212]^and_result204[213]^and_result204[214]^and_result204[215]^and_result204[216]^and_result204[217]^and_result204[218]^and_result204[219]^and_result204[220]^and_result204[221]^and_result204[222]^and_result204[223]^and_result204[224]^and_result204[225]^and_result204[226]^and_result204[227]^and_result204[228]^and_result204[229]^and_result204[230]^and_result204[231]^and_result204[232]^and_result204[233]^and_result204[234]^and_result204[235]^and_result204[236]^and_result204[237]^and_result204[238]^and_result204[239]^and_result204[240]^and_result204[241]^and_result204[242]^and_result204[243]^and_result204[244]^and_result204[245]^and_result204[246]^and_result204[247]^and_result204[248]^and_result204[249]^and_result204[250]^and_result204[251]^and_result204[252]^and_result204[253]^and_result204[254];
assign key[205]=and_result205[0]^and_result205[1]^and_result205[2]^and_result205[3]^and_result205[4]^and_result205[5]^and_result205[6]^and_result205[7]^and_result205[8]^and_result205[9]^and_result205[10]^and_result205[11]^and_result205[12]^and_result205[13]^and_result205[14]^and_result205[15]^and_result205[16]^and_result205[17]^and_result205[18]^and_result205[19]^and_result205[20]^and_result205[21]^and_result205[22]^and_result205[23]^and_result205[24]^and_result205[25]^and_result205[26]^and_result205[27]^and_result205[28]^and_result205[29]^and_result205[30]^and_result205[31]^and_result205[32]^and_result205[33]^and_result205[34]^and_result205[35]^and_result205[36]^and_result205[37]^and_result205[38]^and_result205[39]^and_result205[40]^and_result205[41]^and_result205[42]^and_result205[43]^and_result205[44]^and_result205[45]^and_result205[46]^and_result205[47]^and_result205[48]^and_result205[49]^and_result205[50]^and_result205[51]^and_result205[52]^and_result205[53]^and_result205[54]^and_result205[55]^and_result205[56]^and_result205[57]^and_result205[58]^and_result205[59]^and_result205[60]^and_result205[61]^and_result205[62]^and_result205[63]^and_result205[64]^and_result205[65]^and_result205[66]^and_result205[67]^and_result205[68]^and_result205[69]^and_result205[70]^and_result205[71]^and_result205[72]^and_result205[73]^and_result205[74]^and_result205[75]^and_result205[76]^and_result205[77]^and_result205[78]^and_result205[79]^and_result205[80]^and_result205[81]^and_result205[82]^and_result205[83]^and_result205[84]^and_result205[85]^and_result205[86]^and_result205[87]^and_result205[88]^and_result205[89]^and_result205[90]^and_result205[91]^and_result205[92]^and_result205[93]^and_result205[94]^and_result205[95]^and_result205[96]^and_result205[97]^and_result205[98]^and_result205[99]^and_result205[100]^and_result205[101]^and_result205[102]^and_result205[103]^and_result205[104]^and_result205[105]^and_result205[106]^and_result205[107]^and_result205[108]^and_result205[109]^and_result205[110]^and_result205[111]^and_result205[112]^and_result205[113]^and_result205[114]^and_result205[115]^and_result205[116]^and_result205[117]^and_result205[118]^and_result205[119]^and_result205[120]^and_result205[121]^and_result205[122]^and_result205[123]^and_result205[124]^and_result205[125]^and_result205[126]^and_result205[127]^and_result205[128]^and_result205[129]^and_result205[130]^and_result205[131]^and_result205[132]^and_result205[133]^and_result205[134]^and_result205[135]^and_result205[136]^and_result205[137]^and_result205[138]^and_result205[139]^and_result205[140]^and_result205[141]^and_result205[142]^and_result205[143]^and_result205[144]^and_result205[145]^and_result205[146]^and_result205[147]^and_result205[148]^and_result205[149]^and_result205[150]^and_result205[151]^and_result205[152]^and_result205[153]^and_result205[154]^and_result205[155]^and_result205[156]^and_result205[157]^and_result205[158]^and_result205[159]^and_result205[160]^and_result205[161]^and_result205[162]^and_result205[163]^and_result205[164]^and_result205[165]^and_result205[166]^and_result205[167]^and_result205[168]^and_result205[169]^and_result205[170]^and_result205[171]^and_result205[172]^and_result205[173]^and_result205[174]^and_result205[175]^and_result205[176]^and_result205[177]^and_result205[178]^and_result205[179]^and_result205[180]^and_result205[181]^and_result205[182]^and_result205[183]^and_result205[184]^and_result205[185]^and_result205[186]^and_result205[187]^and_result205[188]^and_result205[189]^and_result205[190]^and_result205[191]^and_result205[192]^and_result205[193]^and_result205[194]^and_result205[195]^and_result205[196]^and_result205[197]^and_result205[198]^and_result205[199]^and_result205[200]^and_result205[201]^and_result205[202]^and_result205[203]^and_result205[204]^and_result205[205]^and_result205[206]^and_result205[207]^and_result205[208]^and_result205[209]^and_result205[210]^and_result205[211]^and_result205[212]^and_result205[213]^and_result205[214]^and_result205[215]^and_result205[216]^and_result205[217]^and_result205[218]^and_result205[219]^and_result205[220]^and_result205[221]^and_result205[222]^and_result205[223]^and_result205[224]^and_result205[225]^and_result205[226]^and_result205[227]^and_result205[228]^and_result205[229]^and_result205[230]^and_result205[231]^and_result205[232]^and_result205[233]^and_result205[234]^and_result205[235]^and_result205[236]^and_result205[237]^and_result205[238]^and_result205[239]^and_result205[240]^and_result205[241]^and_result205[242]^and_result205[243]^and_result205[244]^and_result205[245]^and_result205[246]^and_result205[247]^and_result205[248]^and_result205[249]^and_result205[250]^and_result205[251]^and_result205[252]^and_result205[253]^and_result205[254];
assign key[206]=and_result206[0]^and_result206[1]^and_result206[2]^and_result206[3]^and_result206[4]^and_result206[5]^and_result206[6]^and_result206[7]^and_result206[8]^and_result206[9]^and_result206[10]^and_result206[11]^and_result206[12]^and_result206[13]^and_result206[14]^and_result206[15]^and_result206[16]^and_result206[17]^and_result206[18]^and_result206[19]^and_result206[20]^and_result206[21]^and_result206[22]^and_result206[23]^and_result206[24]^and_result206[25]^and_result206[26]^and_result206[27]^and_result206[28]^and_result206[29]^and_result206[30]^and_result206[31]^and_result206[32]^and_result206[33]^and_result206[34]^and_result206[35]^and_result206[36]^and_result206[37]^and_result206[38]^and_result206[39]^and_result206[40]^and_result206[41]^and_result206[42]^and_result206[43]^and_result206[44]^and_result206[45]^and_result206[46]^and_result206[47]^and_result206[48]^and_result206[49]^and_result206[50]^and_result206[51]^and_result206[52]^and_result206[53]^and_result206[54]^and_result206[55]^and_result206[56]^and_result206[57]^and_result206[58]^and_result206[59]^and_result206[60]^and_result206[61]^and_result206[62]^and_result206[63]^and_result206[64]^and_result206[65]^and_result206[66]^and_result206[67]^and_result206[68]^and_result206[69]^and_result206[70]^and_result206[71]^and_result206[72]^and_result206[73]^and_result206[74]^and_result206[75]^and_result206[76]^and_result206[77]^and_result206[78]^and_result206[79]^and_result206[80]^and_result206[81]^and_result206[82]^and_result206[83]^and_result206[84]^and_result206[85]^and_result206[86]^and_result206[87]^and_result206[88]^and_result206[89]^and_result206[90]^and_result206[91]^and_result206[92]^and_result206[93]^and_result206[94]^and_result206[95]^and_result206[96]^and_result206[97]^and_result206[98]^and_result206[99]^and_result206[100]^and_result206[101]^and_result206[102]^and_result206[103]^and_result206[104]^and_result206[105]^and_result206[106]^and_result206[107]^and_result206[108]^and_result206[109]^and_result206[110]^and_result206[111]^and_result206[112]^and_result206[113]^and_result206[114]^and_result206[115]^and_result206[116]^and_result206[117]^and_result206[118]^and_result206[119]^and_result206[120]^and_result206[121]^and_result206[122]^and_result206[123]^and_result206[124]^and_result206[125]^and_result206[126]^and_result206[127]^and_result206[128]^and_result206[129]^and_result206[130]^and_result206[131]^and_result206[132]^and_result206[133]^and_result206[134]^and_result206[135]^and_result206[136]^and_result206[137]^and_result206[138]^and_result206[139]^and_result206[140]^and_result206[141]^and_result206[142]^and_result206[143]^and_result206[144]^and_result206[145]^and_result206[146]^and_result206[147]^and_result206[148]^and_result206[149]^and_result206[150]^and_result206[151]^and_result206[152]^and_result206[153]^and_result206[154]^and_result206[155]^and_result206[156]^and_result206[157]^and_result206[158]^and_result206[159]^and_result206[160]^and_result206[161]^and_result206[162]^and_result206[163]^and_result206[164]^and_result206[165]^and_result206[166]^and_result206[167]^and_result206[168]^and_result206[169]^and_result206[170]^and_result206[171]^and_result206[172]^and_result206[173]^and_result206[174]^and_result206[175]^and_result206[176]^and_result206[177]^and_result206[178]^and_result206[179]^and_result206[180]^and_result206[181]^and_result206[182]^and_result206[183]^and_result206[184]^and_result206[185]^and_result206[186]^and_result206[187]^and_result206[188]^and_result206[189]^and_result206[190]^and_result206[191]^and_result206[192]^and_result206[193]^and_result206[194]^and_result206[195]^and_result206[196]^and_result206[197]^and_result206[198]^and_result206[199]^and_result206[200]^and_result206[201]^and_result206[202]^and_result206[203]^and_result206[204]^and_result206[205]^and_result206[206]^and_result206[207]^and_result206[208]^and_result206[209]^and_result206[210]^and_result206[211]^and_result206[212]^and_result206[213]^and_result206[214]^and_result206[215]^and_result206[216]^and_result206[217]^and_result206[218]^and_result206[219]^and_result206[220]^and_result206[221]^and_result206[222]^and_result206[223]^and_result206[224]^and_result206[225]^and_result206[226]^and_result206[227]^and_result206[228]^and_result206[229]^and_result206[230]^and_result206[231]^and_result206[232]^and_result206[233]^and_result206[234]^and_result206[235]^and_result206[236]^and_result206[237]^and_result206[238]^and_result206[239]^and_result206[240]^and_result206[241]^and_result206[242]^and_result206[243]^and_result206[244]^and_result206[245]^and_result206[246]^and_result206[247]^and_result206[248]^and_result206[249]^and_result206[250]^and_result206[251]^and_result206[252]^and_result206[253]^and_result206[254];
assign key[207]=and_result207[0]^and_result207[1]^and_result207[2]^and_result207[3]^and_result207[4]^and_result207[5]^and_result207[6]^and_result207[7]^and_result207[8]^and_result207[9]^and_result207[10]^and_result207[11]^and_result207[12]^and_result207[13]^and_result207[14]^and_result207[15]^and_result207[16]^and_result207[17]^and_result207[18]^and_result207[19]^and_result207[20]^and_result207[21]^and_result207[22]^and_result207[23]^and_result207[24]^and_result207[25]^and_result207[26]^and_result207[27]^and_result207[28]^and_result207[29]^and_result207[30]^and_result207[31]^and_result207[32]^and_result207[33]^and_result207[34]^and_result207[35]^and_result207[36]^and_result207[37]^and_result207[38]^and_result207[39]^and_result207[40]^and_result207[41]^and_result207[42]^and_result207[43]^and_result207[44]^and_result207[45]^and_result207[46]^and_result207[47]^and_result207[48]^and_result207[49]^and_result207[50]^and_result207[51]^and_result207[52]^and_result207[53]^and_result207[54]^and_result207[55]^and_result207[56]^and_result207[57]^and_result207[58]^and_result207[59]^and_result207[60]^and_result207[61]^and_result207[62]^and_result207[63]^and_result207[64]^and_result207[65]^and_result207[66]^and_result207[67]^and_result207[68]^and_result207[69]^and_result207[70]^and_result207[71]^and_result207[72]^and_result207[73]^and_result207[74]^and_result207[75]^and_result207[76]^and_result207[77]^and_result207[78]^and_result207[79]^and_result207[80]^and_result207[81]^and_result207[82]^and_result207[83]^and_result207[84]^and_result207[85]^and_result207[86]^and_result207[87]^and_result207[88]^and_result207[89]^and_result207[90]^and_result207[91]^and_result207[92]^and_result207[93]^and_result207[94]^and_result207[95]^and_result207[96]^and_result207[97]^and_result207[98]^and_result207[99]^and_result207[100]^and_result207[101]^and_result207[102]^and_result207[103]^and_result207[104]^and_result207[105]^and_result207[106]^and_result207[107]^and_result207[108]^and_result207[109]^and_result207[110]^and_result207[111]^and_result207[112]^and_result207[113]^and_result207[114]^and_result207[115]^and_result207[116]^and_result207[117]^and_result207[118]^and_result207[119]^and_result207[120]^and_result207[121]^and_result207[122]^and_result207[123]^and_result207[124]^and_result207[125]^and_result207[126]^and_result207[127]^and_result207[128]^and_result207[129]^and_result207[130]^and_result207[131]^and_result207[132]^and_result207[133]^and_result207[134]^and_result207[135]^and_result207[136]^and_result207[137]^and_result207[138]^and_result207[139]^and_result207[140]^and_result207[141]^and_result207[142]^and_result207[143]^and_result207[144]^and_result207[145]^and_result207[146]^and_result207[147]^and_result207[148]^and_result207[149]^and_result207[150]^and_result207[151]^and_result207[152]^and_result207[153]^and_result207[154]^and_result207[155]^and_result207[156]^and_result207[157]^and_result207[158]^and_result207[159]^and_result207[160]^and_result207[161]^and_result207[162]^and_result207[163]^and_result207[164]^and_result207[165]^and_result207[166]^and_result207[167]^and_result207[168]^and_result207[169]^and_result207[170]^and_result207[171]^and_result207[172]^and_result207[173]^and_result207[174]^and_result207[175]^and_result207[176]^and_result207[177]^and_result207[178]^and_result207[179]^and_result207[180]^and_result207[181]^and_result207[182]^and_result207[183]^and_result207[184]^and_result207[185]^and_result207[186]^and_result207[187]^and_result207[188]^and_result207[189]^and_result207[190]^and_result207[191]^and_result207[192]^and_result207[193]^and_result207[194]^and_result207[195]^and_result207[196]^and_result207[197]^and_result207[198]^and_result207[199]^and_result207[200]^and_result207[201]^and_result207[202]^and_result207[203]^and_result207[204]^and_result207[205]^and_result207[206]^and_result207[207]^and_result207[208]^and_result207[209]^and_result207[210]^and_result207[211]^and_result207[212]^and_result207[213]^and_result207[214]^and_result207[215]^and_result207[216]^and_result207[217]^and_result207[218]^and_result207[219]^and_result207[220]^and_result207[221]^and_result207[222]^and_result207[223]^and_result207[224]^and_result207[225]^and_result207[226]^and_result207[227]^and_result207[228]^and_result207[229]^and_result207[230]^and_result207[231]^and_result207[232]^and_result207[233]^and_result207[234]^and_result207[235]^and_result207[236]^and_result207[237]^and_result207[238]^and_result207[239]^and_result207[240]^and_result207[241]^and_result207[242]^and_result207[243]^and_result207[244]^and_result207[245]^and_result207[246]^and_result207[247]^and_result207[248]^and_result207[249]^and_result207[250]^and_result207[251]^and_result207[252]^and_result207[253]^and_result207[254];
assign key[208]=and_result208[0]^and_result208[1]^and_result208[2]^and_result208[3]^and_result208[4]^and_result208[5]^and_result208[6]^and_result208[7]^and_result208[8]^and_result208[9]^and_result208[10]^and_result208[11]^and_result208[12]^and_result208[13]^and_result208[14]^and_result208[15]^and_result208[16]^and_result208[17]^and_result208[18]^and_result208[19]^and_result208[20]^and_result208[21]^and_result208[22]^and_result208[23]^and_result208[24]^and_result208[25]^and_result208[26]^and_result208[27]^and_result208[28]^and_result208[29]^and_result208[30]^and_result208[31]^and_result208[32]^and_result208[33]^and_result208[34]^and_result208[35]^and_result208[36]^and_result208[37]^and_result208[38]^and_result208[39]^and_result208[40]^and_result208[41]^and_result208[42]^and_result208[43]^and_result208[44]^and_result208[45]^and_result208[46]^and_result208[47]^and_result208[48]^and_result208[49]^and_result208[50]^and_result208[51]^and_result208[52]^and_result208[53]^and_result208[54]^and_result208[55]^and_result208[56]^and_result208[57]^and_result208[58]^and_result208[59]^and_result208[60]^and_result208[61]^and_result208[62]^and_result208[63]^and_result208[64]^and_result208[65]^and_result208[66]^and_result208[67]^and_result208[68]^and_result208[69]^and_result208[70]^and_result208[71]^and_result208[72]^and_result208[73]^and_result208[74]^and_result208[75]^and_result208[76]^and_result208[77]^and_result208[78]^and_result208[79]^and_result208[80]^and_result208[81]^and_result208[82]^and_result208[83]^and_result208[84]^and_result208[85]^and_result208[86]^and_result208[87]^and_result208[88]^and_result208[89]^and_result208[90]^and_result208[91]^and_result208[92]^and_result208[93]^and_result208[94]^and_result208[95]^and_result208[96]^and_result208[97]^and_result208[98]^and_result208[99]^and_result208[100]^and_result208[101]^and_result208[102]^and_result208[103]^and_result208[104]^and_result208[105]^and_result208[106]^and_result208[107]^and_result208[108]^and_result208[109]^and_result208[110]^and_result208[111]^and_result208[112]^and_result208[113]^and_result208[114]^and_result208[115]^and_result208[116]^and_result208[117]^and_result208[118]^and_result208[119]^and_result208[120]^and_result208[121]^and_result208[122]^and_result208[123]^and_result208[124]^and_result208[125]^and_result208[126]^and_result208[127]^and_result208[128]^and_result208[129]^and_result208[130]^and_result208[131]^and_result208[132]^and_result208[133]^and_result208[134]^and_result208[135]^and_result208[136]^and_result208[137]^and_result208[138]^and_result208[139]^and_result208[140]^and_result208[141]^and_result208[142]^and_result208[143]^and_result208[144]^and_result208[145]^and_result208[146]^and_result208[147]^and_result208[148]^and_result208[149]^and_result208[150]^and_result208[151]^and_result208[152]^and_result208[153]^and_result208[154]^and_result208[155]^and_result208[156]^and_result208[157]^and_result208[158]^and_result208[159]^and_result208[160]^and_result208[161]^and_result208[162]^and_result208[163]^and_result208[164]^and_result208[165]^and_result208[166]^and_result208[167]^and_result208[168]^and_result208[169]^and_result208[170]^and_result208[171]^and_result208[172]^and_result208[173]^and_result208[174]^and_result208[175]^and_result208[176]^and_result208[177]^and_result208[178]^and_result208[179]^and_result208[180]^and_result208[181]^and_result208[182]^and_result208[183]^and_result208[184]^and_result208[185]^and_result208[186]^and_result208[187]^and_result208[188]^and_result208[189]^and_result208[190]^and_result208[191]^and_result208[192]^and_result208[193]^and_result208[194]^and_result208[195]^and_result208[196]^and_result208[197]^and_result208[198]^and_result208[199]^and_result208[200]^and_result208[201]^and_result208[202]^and_result208[203]^and_result208[204]^and_result208[205]^and_result208[206]^and_result208[207]^and_result208[208]^and_result208[209]^and_result208[210]^and_result208[211]^and_result208[212]^and_result208[213]^and_result208[214]^and_result208[215]^and_result208[216]^and_result208[217]^and_result208[218]^and_result208[219]^and_result208[220]^and_result208[221]^and_result208[222]^and_result208[223]^and_result208[224]^and_result208[225]^and_result208[226]^and_result208[227]^and_result208[228]^and_result208[229]^and_result208[230]^and_result208[231]^and_result208[232]^and_result208[233]^and_result208[234]^and_result208[235]^and_result208[236]^and_result208[237]^and_result208[238]^and_result208[239]^and_result208[240]^and_result208[241]^and_result208[242]^and_result208[243]^and_result208[244]^and_result208[245]^and_result208[246]^and_result208[247]^and_result208[248]^and_result208[249]^and_result208[250]^and_result208[251]^and_result208[252]^and_result208[253]^and_result208[254];
assign key[209]=and_result209[0]^and_result209[1]^and_result209[2]^and_result209[3]^and_result209[4]^and_result209[5]^and_result209[6]^and_result209[7]^and_result209[8]^and_result209[9]^and_result209[10]^and_result209[11]^and_result209[12]^and_result209[13]^and_result209[14]^and_result209[15]^and_result209[16]^and_result209[17]^and_result209[18]^and_result209[19]^and_result209[20]^and_result209[21]^and_result209[22]^and_result209[23]^and_result209[24]^and_result209[25]^and_result209[26]^and_result209[27]^and_result209[28]^and_result209[29]^and_result209[30]^and_result209[31]^and_result209[32]^and_result209[33]^and_result209[34]^and_result209[35]^and_result209[36]^and_result209[37]^and_result209[38]^and_result209[39]^and_result209[40]^and_result209[41]^and_result209[42]^and_result209[43]^and_result209[44]^and_result209[45]^and_result209[46]^and_result209[47]^and_result209[48]^and_result209[49]^and_result209[50]^and_result209[51]^and_result209[52]^and_result209[53]^and_result209[54]^and_result209[55]^and_result209[56]^and_result209[57]^and_result209[58]^and_result209[59]^and_result209[60]^and_result209[61]^and_result209[62]^and_result209[63]^and_result209[64]^and_result209[65]^and_result209[66]^and_result209[67]^and_result209[68]^and_result209[69]^and_result209[70]^and_result209[71]^and_result209[72]^and_result209[73]^and_result209[74]^and_result209[75]^and_result209[76]^and_result209[77]^and_result209[78]^and_result209[79]^and_result209[80]^and_result209[81]^and_result209[82]^and_result209[83]^and_result209[84]^and_result209[85]^and_result209[86]^and_result209[87]^and_result209[88]^and_result209[89]^and_result209[90]^and_result209[91]^and_result209[92]^and_result209[93]^and_result209[94]^and_result209[95]^and_result209[96]^and_result209[97]^and_result209[98]^and_result209[99]^and_result209[100]^and_result209[101]^and_result209[102]^and_result209[103]^and_result209[104]^and_result209[105]^and_result209[106]^and_result209[107]^and_result209[108]^and_result209[109]^and_result209[110]^and_result209[111]^and_result209[112]^and_result209[113]^and_result209[114]^and_result209[115]^and_result209[116]^and_result209[117]^and_result209[118]^and_result209[119]^and_result209[120]^and_result209[121]^and_result209[122]^and_result209[123]^and_result209[124]^and_result209[125]^and_result209[126]^and_result209[127]^and_result209[128]^and_result209[129]^and_result209[130]^and_result209[131]^and_result209[132]^and_result209[133]^and_result209[134]^and_result209[135]^and_result209[136]^and_result209[137]^and_result209[138]^and_result209[139]^and_result209[140]^and_result209[141]^and_result209[142]^and_result209[143]^and_result209[144]^and_result209[145]^and_result209[146]^and_result209[147]^and_result209[148]^and_result209[149]^and_result209[150]^and_result209[151]^and_result209[152]^and_result209[153]^and_result209[154]^and_result209[155]^and_result209[156]^and_result209[157]^and_result209[158]^and_result209[159]^and_result209[160]^and_result209[161]^and_result209[162]^and_result209[163]^and_result209[164]^and_result209[165]^and_result209[166]^and_result209[167]^and_result209[168]^and_result209[169]^and_result209[170]^and_result209[171]^and_result209[172]^and_result209[173]^and_result209[174]^and_result209[175]^and_result209[176]^and_result209[177]^and_result209[178]^and_result209[179]^and_result209[180]^and_result209[181]^and_result209[182]^and_result209[183]^and_result209[184]^and_result209[185]^and_result209[186]^and_result209[187]^and_result209[188]^and_result209[189]^and_result209[190]^and_result209[191]^and_result209[192]^and_result209[193]^and_result209[194]^and_result209[195]^and_result209[196]^and_result209[197]^and_result209[198]^and_result209[199]^and_result209[200]^and_result209[201]^and_result209[202]^and_result209[203]^and_result209[204]^and_result209[205]^and_result209[206]^and_result209[207]^and_result209[208]^and_result209[209]^and_result209[210]^and_result209[211]^and_result209[212]^and_result209[213]^and_result209[214]^and_result209[215]^and_result209[216]^and_result209[217]^and_result209[218]^and_result209[219]^and_result209[220]^and_result209[221]^and_result209[222]^and_result209[223]^and_result209[224]^and_result209[225]^and_result209[226]^and_result209[227]^and_result209[228]^and_result209[229]^and_result209[230]^and_result209[231]^and_result209[232]^and_result209[233]^and_result209[234]^and_result209[235]^and_result209[236]^and_result209[237]^and_result209[238]^and_result209[239]^and_result209[240]^and_result209[241]^and_result209[242]^and_result209[243]^and_result209[244]^and_result209[245]^and_result209[246]^and_result209[247]^and_result209[248]^and_result209[249]^and_result209[250]^and_result209[251]^and_result209[252]^and_result209[253]^and_result209[254];
assign key[210]=and_result210[0]^and_result210[1]^and_result210[2]^and_result210[3]^and_result210[4]^and_result210[5]^and_result210[6]^and_result210[7]^and_result210[8]^and_result210[9]^and_result210[10]^and_result210[11]^and_result210[12]^and_result210[13]^and_result210[14]^and_result210[15]^and_result210[16]^and_result210[17]^and_result210[18]^and_result210[19]^and_result210[20]^and_result210[21]^and_result210[22]^and_result210[23]^and_result210[24]^and_result210[25]^and_result210[26]^and_result210[27]^and_result210[28]^and_result210[29]^and_result210[30]^and_result210[31]^and_result210[32]^and_result210[33]^and_result210[34]^and_result210[35]^and_result210[36]^and_result210[37]^and_result210[38]^and_result210[39]^and_result210[40]^and_result210[41]^and_result210[42]^and_result210[43]^and_result210[44]^and_result210[45]^and_result210[46]^and_result210[47]^and_result210[48]^and_result210[49]^and_result210[50]^and_result210[51]^and_result210[52]^and_result210[53]^and_result210[54]^and_result210[55]^and_result210[56]^and_result210[57]^and_result210[58]^and_result210[59]^and_result210[60]^and_result210[61]^and_result210[62]^and_result210[63]^and_result210[64]^and_result210[65]^and_result210[66]^and_result210[67]^and_result210[68]^and_result210[69]^and_result210[70]^and_result210[71]^and_result210[72]^and_result210[73]^and_result210[74]^and_result210[75]^and_result210[76]^and_result210[77]^and_result210[78]^and_result210[79]^and_result210[80]^and_result210[81]^and_result210[82]^and_result210[83]^and_result210[84]^and_result210[85]^and_result210[86]^and_result210[87]^and_result210[88]^and_result210[89]^and_result210[90]^and_result210[91]^and_result210[92]^and_result210[93]^and_result210[94]^and_result210[95]^and_result210[96]^and_result210[97]^and_result210[98]^and_result210[99]^and_result210[100]^and_result210[101]^and_result210[102]^and_result210[103]^and_result210[104]^and_result210[105]^and_result210[106]^and_result210[107]^and_result210[108]^and_result210[109]^and_result210[110]^and_result210[111]^and_result210[112]^and_result210[113]^and_result210[114]^and_result210[115]^and_result210[116]^and_result210[117]^and_result210[118]^and_result210[119]^and_result210[120]^and_result210[121]^and_result210[122]^and_result210[123]^and_result210[124]^and_result210[125]^and_result210[126]^and_result210[127]^and_result210[128]^and_result210[129]^and_result210[130]^and_result210[131]^and_result210[132]^and_result210[133]^and_result210[134]^and_result210[135]^and_result210[136]^and_result210[137]^and_result210[138]^and_result210[139]^and_result210[140]^and_result210[141]^and_result210[142]^and_result210[143]^and_result210[144]^and_result210[145]^and_result210[146]^and_result210[147]^and_result210[148]^and_result210[149]^and_result210[150]^and_result210[151]^and_result210[152]^and_result210[153]^and_result210[154]^and_result210[155]^and_result210[156]^and_result210[157]^and_result210[158]^and_result210[159]^and_result210[160]^and_result210[161]^and_result210[162]^and_result210[163]^and_result210[164]^and_result210[165]^and_result210[166]^and_result210[167]^and_result210[168]^and_result210[169]^and_result210[170]^and_result210[171]^and_result210[172]^and_result210[173]^and_result210[174]^and_result210[175]^and_result210[176]^and_result210[177]^and_result210[178]^and_result210[179]^and_result210[180]^and_result210[181]^and_result210[182]^and_result210[183]^and_result210[184]^and_result210[185]^and_result210[186]^and_result210[187]^and_result210[188]^and_result210[189]^and_result210[190]^and_result210[191]^and_result210[192]^and_result210[193]^and_result210[194]^and_result210[195]^and_result210[196]^and_result210[197]^and_result210[198]^and_result210[199]^and_result210[200]^and_result210[201]^and_result210[202]^and_result210[203]^and_result210[204]^and_result210[205]^and_result210[206]^and_result210[207]^and_result210[208]^and_result210[209]^and_result210[210]^and_result210[211]^and_result210[212]^and_result210[213]^and_result210[214]^and_result210[215]^and_result210[216]^and_result210[217]^and_result210[218]^and_result210[219]^and_result210[220]^and_result210[221]^and_result210[222]^and_result210[223]^and_result210[224]^and_result210[225]^and_result210[226]^and_result210[227]^and_result210[228]^and_result210[229]^and_result210[230]^and_result210[231]^and_result210[232]^and_result210[233]^and_result210[234]^and_result210[235]^and_result210[236]^and_result210[237]^and_result210[238]^and_result210[239]^and_result210[240]^and_result210[241]^and_result210[242]^and_result210[243]^and_result210[244]^and_result210[245]^and_result210[246]^and_result210[247]^and_result210[248]^and_result210[249]^and_result210[250]^and_result210[251]^and_result210[252]^and_result210[253]^and_result210[254];
assign key[211]=and_result211[0]^and_result211[1]^and_result211[2]^and_result211[3]^and_result211[4]^and_result211[5]^and_result211[6]^and_result211[7]^and_result211[8]^and_result211[9]^and_result211[10]^and_result211[11]^and_result211[12]^and_result211[13]^and_result211[14]^and_result211[15]^and_result211[16]^and_result211[17]^and_result211[18]^and_result211[19]^and_result211[20]^and_result211[21]^and_result211[22]^and_result211[23]^and_result211[24]^and_result211[25]^and_result211[26]^and_result211[27]^and_result211[28]^and_result211[29]^and_result211[30]^and_result211[31]^and_result211[32]^and_result211[33]^and_result211[34]^and_result211[35]^and_result211[36]^and_result211[37]^and_result211[38]^and_result211[39]^and_result211[40]^and_result211[41]^and_result211[42]^and_result211[43]^and_result211[44]^and_result211[45]^and_result211[46]^and_result211[47]^and_result211[48]^and_result211[49]^and_result211[50]^and_result211[51]^and_result211[52]^and_result211[53]^and_result211[54]^and_result211[55]^and_result211[56]^and_result211[57]^and_result211[58]^and_result211[59]^and_result211[60]^and_result211[61]^and_result211[62]^and_result211[63]^and_result211[64]^and_result211[65]^and_result211[66]^and_result211[67]^and_result211[68]^and_result211[69]^and_result211[70]^and_result211[71]^and_result211[72]^and_result211[73]^and_result211[74]^and_result211[75]^and_result211[76]^and_result211[77]^and_result211[78]^and_result211[79]^and_result211[80]^and_result211[81]^and_result211[82]^and_result211[83]^and_result211[84]^and_result211[85]^and_result211[86]^and_result211[87]^and_result211[88]^and_result211[89]^and_result211[90]^and_result211[91]^and_result211[92]^and_result211[93]^and_result211[94]^and_result211[95]^and_result211[96]^and_result211[97]^and_result211[98]^and_result211[99]^and_result211[100]^and_result211[101]^and_result211[102]^and_result211[103]^and_result211[104]^and_result211[105]^and_result211[106]^and_result211[107]^and_result211[108]^and_result211[109]^and_result211[110]^and_result211[111]^and_result211[112]^and_result211[113]^and_result211[114]^and_result211[115]^and_result211[116]^and_result211[117]^and_result211[118]^and_result211[119]^and_result211[120]^and_result211[121]^and_result211[122]^and_result211[123]^and_result211[124]^and_result211[125]^and_result211[126]^and_result211[127]^and_result211[128]^and_result211[129]^and_result211[130]^and_result211[131]^and_result211[132]^and_result211[133]^and_result211[134]^and_result211[135]^and_result211[136]^and_result211[137]^and_result211[138]^and_result211[139]^and_result211[140]^and_result211[141]^and_result211[142]^and_result211[143]^and_result211[144]^and_result211[145]^and_result211[146]^and_result211[147]^and_result211[148]^and_result211[149]^and_result211[150]^and_result211[151]^and_result211[152]^and_result211[153]^and_result211[154]^and_result211[155]^and_result211[156]^and_result211[157]^and_result211[158]^and_result211[159]^and_result211[160]^and_result211[161]^and_result211[162]^and_result211[163]^and_result211[164]^and_result211[165]^and_result211[166]^and_result211[167]^and_result211[168]^and_result211[169]^and_result211[170]^and_result211[171]^and_result211[172]^and_result211[173]^and_result211[174]^and_result211[175]^and_result211[176]^and_result211[177]^and_result211[178]^and_result211[179]^and_result211[180]^and_result211[181]^and_result211[182]^and_result211[183]^and_result211[184]^and_result211[185]^and_result211[186]^and_result211[187]^and_result211[188]^and_result211[189]^and_result211[190]^and_result211[191]^and_result211[192]^and_result211[193]^and_result211[194]^and_result211[195]^and_result211[196]^and_result211[197]^and_result211[198]^and_result211[199]^and_result211[200]^and_result211[201]^and_result211[202]^and_result211[203]^and_result211[204]^and_result211[205]^and_result211[206]^and_result211[207]^and_result211[208]^and_result211[209]^and_result211[210]^and_result211[211]^and_result211[212]^and_result211[213]^and_result211[214]^and_result211[215]^and_result211[216]^and_result211[217]^and_result211[218]^and_result211[219]^and_result211[220]^and_result211[221]^and_result211[222]^and_result211[223]^and_result211[224]^and_result211[225]^and_result211[226]^and_result211[227]^and_result211[228]^and_result211[229]^and_result211[230]^and_result211[231]^and_result211[232]^and_result211[233]^and_result211[234]^and_result211[235]^and_result211[236]^and_result211[237]^and_result211[238]^and_result211[239]^and_result211[240]^and_result211[241]^and_result211[242]^and_result211[243]^and_result211[244]^and_result211[245]^and_result211[246]^and_result211[247]^and_result211[248]^and_result211[249]^and_result211[250]^and_result211[251]^and_result211[252]^and_result211[253]^and_result211[254];
assign key[212]=and_result212[0]^and_result212[1]^and_result212[2]^and_result212[3]^and_result212[4]^and_result212[5]^and_result212[6]^and_result212[7]^and_result212[8]^and_result212[9]^and_result212[10]^and_result212[11]^and_result212[12]^and_result212[13]^and_result212[14]^and_result212[15]^and_result212[16]^and_result212[17]^and_result212[18]^and_result212[19]^and_result212[20]^and_result212[21]^and_result212[22]^and_result212[23]^and_result212[24]^and_result212[25]^and_result212[26]^and_result212[27]^and_result212[28]^and_result212[29]^and_result212[30]^and_result212[31]^and_result212[32]^and_result212[33]^and_result212[34]^and_result212[35]^and_result212[36]^and_result212[37]^and_result212[38]^and_result212[39]^and_result212[40]^and_result212[41]^and_result212[42]^and_result212[43]^and_result212[44]^and_result212[45]^and_result212[46]^and_result212[47]^and_result212[48]^and_result212[49]^and_result212[50]^and_result212[51]^and_result212[52]^and_result212[53]^and_result212[54]^and_result212[55]^and_result212[56]^and_result212[57]^and_result212[58]^and_result212[59]^and_result212[60]^and_result212[61]^and_result212[62]^and_result212[63]^and_result212[64]^and_result212[65]^and_result212[66]^and_result212[67]^and_result212[68]^and_result212[69]^and_result212[70]^and_result212[71]^and_result212[72]^and_result212[73]^and_result212[74]^and_result212[75]^and_result212[76]^and_result212[77]^and_result212[78]^and_result212[79]^and_result212[80]^and_result212[81]^and_result212[82]^and_result212[83]^and_result212[84]^and_result212[85]^and_result212[86]^and_result212[87]^and_result212[88]^and_result212[89]^and_result212[90]^and_result212[91]^and_result212[92]^and_result212[93]^and_result212[94]^and_result212[95]^and_result212[96]^and_result212[97]^and_result212[98]^and_result212[99]^and_result212[100]^and_result212[101]^and_result212[102]^and_result212[103]^and_result212[104]^and_result212[105]^and_result212[106]^and_result212[107]^and_result212[108]^and_result212[109]^and_result212[110]^and_result212[111]^and_result212[112]^and_result212[113]^and_result212[114]^and_result212[115]^and_result212[116]^and_result212[117]^and_result212[118]^and_result212[119]^and_result212[120]^and_result212[121]^and_result212[122]^and_result212[123]^and_result212[124]^and_result212[125]^and_result212[126]^and_result212[127]^and_result212[128]^and_result212[129]^and_result212[130]^and_result212[131]^and_result212[132]^and_result212[133]^and_result212[134]^and_result212[135]^and_result212[136]^and_result212[137]^and_result212[138]^and_result212[139]^and_result212[140]^and_result212[141]^and_result212[142]^and_result212[143]^and_result212[144]^and_result212[145]^and_result212[146]^and_result212[147]^and_result212[148]^and_result212[149]^and_result212[150]^and_result212[151]^and_result212[152]^and_result212[153]^and_result212[154]^and_result212[155]^and_result212[156]^and_result212[157]^and_result212[158]^and_result212[159]^and_result212[160]^and_result212[161]^and_result212[162]^and_result212[163]^and_result212[164]^and_result212[165]^and_result212[166]^and_result212[167]^and_result212[168]^and_result212[169]^and_result212[170]^and_result212[171]^and_result212[172]^and_result212[173]^and_result212[174]^and_result212[175]^and_result212[176]^and_result212[177]^and_result212[178]^and_result212[179]^and_result212[180]^and_result212[181]^and_result212[182]^and_result212[183]^and_result212[184]^and_result212[185]^and_result212[186]^and_result212[187]^and_result212[188]^and_result212[189]^and_result212[190]^and_result212[191]^and_result212[192]^and_result212[193]^and_result212[194]^and_result212[195]^and_result212[196]^and_result212[197]^and_result212[198]^and_result212[199]^and_result212[200]^and_result212[201]^and_result212[202]^and_result212[203]^and_result212[204]^and_result212[205]^and_result212[206]^and_result212[207]^and_result212[208]^and_result212[209]^and_result212[210]^and_result212[211]^and_result212[212]^and_result212[213]^and_result212[214]^and_result212[215]^and_result212[216]^and_result212[217]^and_result212[218]^and_result212[219]^and_result212[220]^and_result212[221]^and_result212[222]^and_result212[223]^and_result212[224]^and_result212[225]^and_result212[226]^and_result212[227]^and_result212[228]^and_result212[229]^and_result212[230]^and_result212[231]^and_result212[232]^and_result212[233]^and_result212[234]^and_result212[235]^and_result212[236]^and_result212[237]^and_result212[238]^and_result212[239]^and_result212[240]^and_result212[241]^and_result212[242]^and_result212[243]^and_result212[244]^and_result212[245]^and_result212[246]^and_result212[247]^and_result212[248]^and_result212[249]^and_result212[250]^and_result212[251]^and_result212[252]^and_result212[253]^and_result212[254];
assign key[213]=and_result213[0]^and_result213[1]^and_result213[2]^and_result213[3]^and_result213[4]^and_result213[5]^and_result213[6]^and_result213[7]^and_result213[8]^and_result213[9]^and_result213[10]^and_result213[11]^and_result213[12]^and_result213[13]^and_result213[14]^and_result213[15]^and_result213[16]^and_result213[17]^and_result213[18]^and_result213[19]^and_result213[20]^and_result213[21]^and_result213[22]^and_result213[23]^and_result213[24]^and_result213[25]^and_result213[26]^and_result213[27]^and_result213[28]^and_result213[29]^and_result213[30]^and_result213[31]^and_result213[32]^and_result213[33]^and_result213[34]^and_result213[35]^and_result213[36]^and_result213[37]^and_result213[38]^and_result213[39]^and_result213[40]^and_result213[41]^and_result213[42]^and_result213[43]^and_result213[44]^and_result213[45]^and_result213[46]^and_result213[47]^and_result213[48]^and_result213[49]^and_result213[50]^and_result213[51]^and_result213[52]^and_result213[53]^and_result213[54]^and_result213[55]^and_result213[56]^and_result213[57]^and_result213[58]^and_result213[59]^and_result213[60]^and_result213[61]^and_result213[62]^and_result213[63]^and_result213[64]^and_result213[65]^and_result213[66]^and_result213[67]^and_result213[68]^and_result213[69]^and_result213[70]^and_result213[71]^and_result213[72]^and_result213[73]^and_result213[74]^and_result213[75]^and_result213[76]^and_result213[77]^and_result213[78]^and_result213[79]^and_result213[80]^and_result213[81]^and_result213[82]^and_result213[83]^and_result213[84]^and_result213[85]^and_result213[86]^and_result213[87]^and_result213[88]^and_result213[89]^and_result213[90]^and_result213[91]^and_result213[92]^and_result213[93]^and_result213[94]^and_result213[95]^and_result213[96]^and_result213[97]^and_result213[98]^and_result213[99]^and_result213[100]^and_result213[101]^and_result213[102]^and_result213[103]^and_result213[104]^and_result213[105]^and_result213[106]^and_result213[107]^and_result213[108]^and_result213[109]^and_result213[110]^and_result213[111]^and_result213[112]^and_result213[113]^and_result213[114]^and_result213[115]^and_result213[116]^and_result213[117]^and_result213[118]^and_result213[119]^and_result213[120]^and_result213[121]^and_result213[122]^and_result213[123]^and_result213[124]^and_result213[125]^and_result213[126]^and_result213[127]^and_result213[128]^and_result213[129]^and_result213[130]^and_result213[131]^and_result213[132]^and_result213[133]^and_result213[134]^and_result213[135]^and_result213[136]^and_result213[137]^and_result213[138]^and_result213[139]^and_result213[140]^and_result213[141]^and_result213[142]^and_result213[143]^and_result213[144]^and_result213[145]^and_result213[146]^and_result213[147]^and_result213[148]^and_result213[149]^and_result213[150]^and_result213[151]^and_result213[152]^and_result213[153]^and_result213[154]^and_result213[155]^and_result213[156]^and_result213[157]^and_result213[158]^and_result213[159]^and_result213[160]^and_result213[161]^and_result213[162]^and_result213[163]^and_result213[164]^and_result213[165]^and_result213[166]^and_result213[167]^and_result213[168]^and_result213[169]^and_result213[170]^and_result213[171]^and_result213[172]^and_result213[173]^and_result213[174]^and_result213[175]^and_result213[176]^and_result213[177]^and_result213[178]^and_result213[179]^and_result213[180]^and_result213[181]^and_result213[182]^and_result213[183]^and_result213[184]^and_result213[185]^and_result213[186]^and_result213[187]^and_result213[188]^and_result213[189]^and_result213[190]^and_result213[191]^and_result213[192]^and_result213[193]^and_result213[194]^and_result213[195]^and_result213[196]^and_result213[197]^and_result213[198]^and_result213[199]^and_result213[200]^and_result213[201]^and_result213[202]^and_result213[203]^and_result213[204]^and_result213[205]^and_result213[206]^and_result213[207]^and_result213[208]^and_result213[209]^and_result213[210]^and_result213[211]^and_result213[212]^and_result213[213]^and_result213[214]^and_result213[215]^and_result213[216]^and_result213[217]^and_result213[218]^and_result213[219]^and_result213[220]^and_result213[221]^and_result213[222]^and_result213[223]^and_result213[224]^and_result213[225]^and_result213[226]^and_result213[227]^and_result213[228]^and_result213[229]^and_result213[230]^and_result213[231]^and_result213[232]^and_result213[233]^and_result213[234]^and_result213[235]^and_result213[236]^and_result213[237]^and_result213[238]^and_result213[239]^and_result213[240]^and_result213[241]^and_result213[242]^and_result213[243]^and_result213[244]^and_result213[245]^and_result213[246]^and_result213[247]^and_result213[248]^and_result213[249]^and_result213[250]^and_result213[251]^and_result213[252]^and_result213[253]^and_result213[254];
assign key[214]=and_result214[0]^and_result214[1]^and_result214[2]^and_result214[3]^and_result214[4]^and_result214[5]^and_result214[6]^and_result214[7]^and_result214[8]^and_result214[9]^and_result214[10]^and_result214[11]^and_result214[12]^and_result214[13]^and_result214[14]^and_result214[15]^and_result214[16]^and_result214[17]^and_result214[18]^and_result214[19]^and_result214[20]^and_result214[21]^and_result214[22]^and_result214[23]^and_result214[24]^and_result214[25]^and_result214[26]^and_result214[27]^and_result214[28]^and_result214[29]^and_result214[30]^and_result214[31]^and_result214[32]^and_result214[33]^and_result214[34]^and_result214[35]^and_result214[36]^and_result214[37]^and_result214[38]^and_result214[39]^and_result214[40]^and_result214[41]^and_result214[42]^and_result214[43]^and_result214[44]^and_result214[45]^and_result214[46]^and_result214[47]^and_result214[48]^and_result214[49]^and_result214[50]^and_result214[51]^and_result214[52]^and_result214[53]^and_result214[54]^and_result214[55]^and_result214[56]^and_result214[57]^and_result214[58]^and_result214[59]^and_result214[60]^and_result214[61]^and_result214[62]^and_result214[63]^and_result214[64]^and_result214[65]^and_result214[66]^and_result214[67]^and_result214[68]^and_result214[69]^and_result214[70]^and_result214[71]^and_result214[72]^and_result214[73]^and_result214[74]^and_result214[75]^and_result214[76]^and_result214[77]^and_result214[78]^and_result214[79]^and_result214[80]^and_result214[81]^and_result214[82]^and_result214[83]^and_result214[84]^and_result214[85]^and_result214[86]^and_result214[87]^and_result214[88]^and_result214[89]^and_result214[90]^and_result214[91]^and_result214[92]^and_result214[93]^and_result214[94]^and_result214[95]^and_result214[96]^and_result214[97]^and_result214[98]^and_result214[99]^and_result214[100]^and_result214[101]^and_result214[102]^and_result214[103]^and_result214[104]^and_result214[105]^and_result214[106]^and_result214[107]^and_result214[108]^and_result214[109]^and_result214[110]^and_result214[111]^and_result214[112]^and_result214[113]^and_result214[114]^and_result214[115]^and_result214[116]^and_result214[117]^and_result214[118]^and_result214[119]^and_result214[120]^and_result214[121]^and_result214[122]^and_result214[123]^and_result214[124]^and_result214[125]^and_result214[126]^and_result214[127]^and_result214[128]^and_result214[129]^and_result214[130]^and_result214[131]^and_result214[132]^and_result214[133]^and_result214[134]^and_result214[135]^and_result214[136]^and_result214[137]^and_result214[138]^and_result214[139]^and_result214[140]^and_result214[141]^and_result214[142]^and_result214[143]^and_result214[144]^and_result214[145]^and_result214[146]^and_result214[147]^and_result214[148]^and_result214[149]^and_result214[150]^and_result214[151]^and_result214[152]^and_result214[153]^and_result214[154]^and_result214[155]^and_result214[156]^and_result214[157]^and_result214[158]^and_result214[159]^and_result214[160]^and_result214[161]^and_result214[162]^and_result214[163]^and_result214[164]^and_result214[165]^and_result214[166]^and_result214[167]^and_result214[168]^and_result214[169]^and_result214[170]^and_result214[171]^and_result214[172]^and_result214[173]^and_result214[174]^and_result214[175]^and_result214[176]^and_result214[177]^and_result214[178]^and_result214[179]^and_result214[180]^and_result214[181]^and_result214[182]^and_result214[183]^and_result214[184]^and_result214[185]^and_result214[186]^and_result214[187]^and_result214[188]^and_result214[189]^and_result214[190]^and_result214[191]^and_result214[192]^and_result214[193]^and_result214[194]^and_result214[195]^and_result214[196]^and_result214[197]^and_result214[198]^and_result214[199]^and_result214[200]^and_result214[201]^and_result214[202]^and_result214[203]^and_result214[204]^and_result214[205]^and_result214[206]^and_result214[207]^and_result214[208]^and_result214[209]^and_result214[210]^and_result214[211]^and_result214[212]^and_result214[213]^and_result214[214]^and_result214[215]^and_result214[216]^and_result214[217]^and_result214[218]^and_result214[219]^and_result214[220]^and_result214[221]^and_result214[222]^and_result214[223]^and_result214[224]^and_result214[225]^and_result214[226]^and_result214[227]^and_result214[228]^and_result214[229]^and_result214[230]^and_result214[231]^and_result214[232]^and_result214[233]^and_result214[234]^and_result214[235]^and_result214[236]^and_result214[237]^and_result214[238]^and_result214[239]^and_result214[240]^and_result214[241]^and_result214[242]^and_result214[243]^and_result214[244]^and_result214[245]^and_result214[246]^and_result214[247]^and_result214[248]^and_result214[249]^and_result214[250]^and_result214[251]^and_result214[252]^and_result214[253]^and_result214[254];
assign key[215]=and_result215[0]^and_result215[1]^and_result215[2]^and_result215[3]^and_result215[4]^and_result215[5]^and_result215[6]^and_result215[7]^and_result215[8]^and_result215[9]^and_result215[10]^and_result215[11]^and_result215[12]^and_result215[13]^and_result215[14]^and_result215[15]^and_result215[16]^and_result215[17]^and_result215[18]^and_result215[19]^and_result215[20]^and_result215[21]^and_result215[22]^and_result215[23]^and_result215[24]^and_result215[25]^and_result215[26]^and_result215[27]^and_result215[28]^and_result215[29]^and_result215[30]^and_result215[31]^and_result215[32]^and_result215[33]^and_result215[34]^and_result215[35]^and_result215[36]^and_result215[37]^and_result215[38]^and_result215[39]^and_result215[40]^and_result215[41]^and_result215[42]^and_result215[43]^and_result215[44]^and_result215[45]^and_result215[46]^and_result215[47]^and_result215[48]^and_result215[49]^and_result215[50]^and_result215[51]^and_result215[52]^and_result215[53]^and_result215[54]^and_result215[55]^and_result215[56]^and_result215[57]^and_result215[58]^and_result215[59]^and_result215[60]^and_result215[61]^and_result215[62]^and_result215[63]^and_result215[64]^and_result215[65]^and_result215[66]^and_result215[67]^and_result215[68]^and_result215[69]^and_result215[70]^and_result215[71]^and_result215[72]^and_result215[73]^and_result215[74]^and_result215[75]^and_result215[76]^and_result215[77]^and_result215[78]^and_result215[79]^and_result215[80]^and_result215[81]^and_result215[82]^and_result215[83]^and_result215[84]^and_result215[85]^and_result215[86]^and_result215[87]^and_result215[88]^and_result215[89]^and_result215[90]^and_result215[91]^and_result215[92]^and_result215[93]^and_result215[94]^and_result215[95]^and_result215[96]^and_result215[97]^and_result215[98]^and_result215[99]^and_result215[100]^and_result215[101]^and_result215[102]^and_result215[103]^and_result215[104]^and_result215[105]^and_result215[106]^and_result215[107]^and_result215[108]^and_result215[109]^and_result215[110]^and_result215[111]^and_result215[112]^and_result215[113]^and_result215[114]^and_result215[115]^and_result215[116]^and_result215[117]^and_result215[118]^and_result215[119]^and_result215[120]^and_result215[121]^and_result215[122]^and_result215[123]^and_result215[124]^and_result215[125]^and_result215[126]^and_result215[127]^and_result215[128]^and_result215[129]^and_result215[130]^and_result215[131]^and_result215[132]^and_result215[133]^and_result215[134]^and_result215[135]^and_result215[136]^and_result215[137]^and_result215[138]^and_result215[139]^and_result215[140]^and_result215[141]^and_result215[142]^and_result215[143]^and_result215[144]^and_result215[145]^and_result215[146]^and_result215[147]^and_result215[148]^and_result215[149]^and_result215[150]^and_result215[151]^and_result215[152]^and_result215[153]^and_result215[154]^and_result215[155]^and_result215[156]^and_result215[157]^and_result215[158]^and_result215[159]^and_result215[160]^and_result215[161]^and_result215[162]^and_result215[163]^and_result215[164]^and_result215[165]^and_result215[166]^and_result215[167]^and_result215[168]^and_result215[169]^and_result215[170]^and_result215[171]^and_result215[172]^and_result215[173]^and_result215[174]^and_result215[175]^and_result215[176]^and_result215[177]^and_result215[178]^and_result215[179]^and_result215[180]^and_result215[181]^and_result215[182]^and_result215[183]^and_result215[184]^and_result215[185]^and_result215[186]^and_result215[187]^and_result215[188]^and_result215[189]^and_result215[190]^and_result215[191]^and_result215[192]^and_result215[193]^and_result215[194]^and_result215[195]^and_result215[196]^and_result215[197]^and_result215[198]^and_result215[199]^and_result215[200]^and_result215[201]^and_result215[202]^and_result215[203]^and_result215[204]^and_result215[205]^and_result215[206]^and_result215[207]^and_result215[208]^and_result215[209]^and_result215[210]^and_result215[211]^and_result215[212]^and_result215[213]^and_result215[214]^and_result215[215]^and_result215[216]^and_result215[217]^and_result215[218]^and_result215[219]^and_result215[220]^and_result215[221]^and_result215[222]^and_result215[223]^and_result215[224]^and_result215[225]^and_result215[226]^and_result215[227]^and_result215[228]^and_result215[229]^and_result215[230]^and_result215[231]^and_result215[232]^and_result215[233]^and_result215[234]^and_result215[235]^and_result215[236]^and_result215[237]^and_result215[238]^and_result215[239]^and_result215[240]^and_result215[241]^and_result215[242]^and_result215[243]^and_result215[244]^and_result215[245]^and_result215[246]^and_result215[247]^and_result215[248]^and_result215[249]^and_result215[250]^and_result215[251]^and_result215[252]^and_result215[253]^and_result215[254];
assign key[216]=and_result216[0]^and_result216[1]^and_result216[2]^and_result216[3]^and_result216[4]^and_result216[5]^and_result216[6]^and_result216[7]^and_result216[8]^and_result216[9]^and_result216[10]^and_result216[11]^and_result216[12]^and_result216[13]^and_result216[14]^and_result216[15]^and_result216[16]^and_result216[17]^and_result216[18]^and_result216[19]^and_result216[20]^and_result216[21]^and_result216[22]^and_result216[23]^and_result216[24]^and_result216[25]^and_result216[26]^and_result216[27]^and_result216[28]^and_result216[29]^and_result216[30]^and_result216[31]^and_result216[32]^and_result216[33]^and_result216[34]^and_result216[35]^and_result216[36]^and_result216[37]^and_result216[38]^and_result216[39]^and_result216[40]^and_result216[41]^and_result216[42]^and_result216[43]^and_result216[44]^and_result216[45]^and_result216[46]^and_result216[47]^and_result216[48]^and_result216[49]^and_result216[50]^and_result216[51]^and_result216[52]^and_result216[53]^and_result216[54]^and_result216[55]^and_result216[56]^and_result216[57]^and_result216[58]^and_result216[59]^and_result216[60]^and_result216[61]^and_result216[62]^and_result216[63]^and_result216[64]^and_result216[65]^and_result216[66]^and_result216[67]^and_result216[68]^and_result216[69]^and_result216[70]^and_result216[71]^and_result216[72]^and_result216[73]^and_result216[74]^and_result216[75]^and_result216[76]^and_result216[77]^and_result216[78]^and_result216[79]^and_result216[80]^and_result216[81]^and_result216[82]^and_result216[83]^and_result216[84]^and_result216[85]^and_result216[86]^and_result216[87]^and_result216[88]^and_result216[89]^and_result216[90]^and_result216[91]^and_result216[92]^and_result216[93]^and_result216[94]^and_result216[95]^and_result216[96]^and_result216[97]^and_result216[98]^and_result216[99]^and_result216[100]^and_result216[101]^and_result216[102]^and_result216[103]^and_result216[104]^and_result216[105]^and_result216[106]^and_result216[107]^and_result216[108]^and_result216[109]^and_result216[110]^and_result216[111]^and_result216[112]^and_result216[113]^and_result216[114]^and_result216[115]^and_result216[116]^and_result216[117]^and_result216[118]^and_result216[119]^and_result216[120]^and_result216[121]^and_result216[122]^and_result216[123]^and_result216[124]^and_result216[125]^and_result216[126]^and_result216[127]^and_result216[128]^and_result216[129]^and_result216[130]^and_result216[131]^and_result216[132]^and_result216[133]^and_result216[134]^and_result216[135]^and_result216[136]^and_result216[137]^and_result216[138]^and_result216[139]^and_result216[140]^and_result216[141]^and_result216[142]^and_result216[143]^and_result216[144]^and_result216[145]^and_result216[146]^and_result216[147]^and_result216[148]^and_result216[149]^and_result216[150]^and_result216[151]^and_result216[152]^and_result216[153]^and_result216[154]^and_result216[155]^and_result216[156]^and_result216[157]^and_result216[158]^and_result216[159]^and_result216[160]^and_result216[161]^and_result216[162]^and_result216[163]^and_result216[164]^and_result216[165]^and_result216[166]^and_result216[167]^and_result216[168]^and_result216[169]^and_result216[170]^and_result216[171]^and_result216[172]^and_result216[173]^and_result216[174]^and_result216[175]^and_result216[176]^and_result216[177]^and_result216[178]^and_result216[179]^and_result216[180]^and_result216[181]^and_result216[182]^and_result216[183]^and_result216[184]^and_result216[185]^and_result216[186]^and_result216[187]^and_result216[188]^and_result216[189]^and_result216[190]^and_result216[191]^and_result216[192]^and_result216[193]^and_result216[194]^and_result216[195]^and_result216[196]^and_result216[197]^and_result216[198]^and_result216[199]^and_result216[200]^and_result216[201]^and_result216[202]^and_result216[203]^and_result216[204]^and_result216[205]^and_result216[206]^and_result216[207]^and_result216[208]^and_result216[209]^and_result216[210]^and_result216[211]^and_result216[212]^and_result216[213]^and_result216[214]^and_result216[215]^and_result216[216]^and_result216[217]^and_result216[218]^and_result216[219]^and_result216[220]^and_result216[221]^and_result216[222]^and_result216[223]^and_result216[224]^and_result216[225]^and_result216[226]^and_result216[227]^and_result216[228]^and_result216[229]^and_result216[230]^and_result216[231]^and_result216[232]^and_result216[233]^and_result216[234]^and_result216[235]^and_result216[236]^and_result216[237]^and_result216[238]^and_result216[239]^and_result216[240]^and_result216[241]^and_result216[242]^and_result216[243]^and_result216[244]^and_result216[245]^and_result216[246]^and_result216[247]^and_result216[248]^and_result216[249]^and_result216[250]^and_result216[251]^and_result216[252]^and_result216[253]^and_result216[254];
assign key[217]=and_result217[0]^and_result217[1]^and_result217[2]^and_result217[3]^and_result217[4]^and_result217[5]^and_result217[6]^and_result217[7]^and_result217[8]^and_result217[9]^and_result217[10]^and_result217[11]^and_result217[12]^and_result217[13]^and_result217[14]^and_result217[15]^and_result217[16]^and_result217[17]^and_result217[18]^and_result217[19]^and_result217[20]^and_result217[21]^and_result217[22]^and_result217[23]^and_result217[24]^and_result217[25]^and_result217[26]^and_result217[27]^and_result217[28]^and_result217[29]^and_result217[30]^and_result217[31]^and_result217[32]^and_result217[33]^and_result217[34]^and_result217[35]^and_result217[36]^and_result217[37]^and_result217[38]^and_result217[39]^and_result217[40]^and_result217[41]^and_result217[42]^and_result217[43]^and_result217[44]^and_result217[45]^and_result217[46]^and_result217[47]^and_result217[48]^and_result217[49]^and_result217[50]^and_result217[51]^and_result217[52]^and_result217[53]^and_result217[54]^and_result217[55]^and_result217[56]^and_result217[57]^and_result217[58]^and_result217[59]^and_result217[60]^and_result217[61]^and_result217[62]^and_result217[63]^and_result217[64]^and_result217[65]^and_result217[66]^and_result217[67]^and_result217[68]^and_result217[69]^and_result217[70]^and_result217[71]^and_result217[72]^and_result217[73]^and_result217[74]^and_result217[75]^and_result217[76]^and_result217[77]^and_result217[78]^and_result217[79]^and_result217[80]^and_result217[81]^and_result217[82]^and_result217[83]^and_result217[84]^and_result217[85]^and_result217[86]^and_result217[87]^and_result217[88]^and_result217[89]^and_result217[90]^and_result217[91]^and_result217[92]^and_result217[93]^and_result217[94]^and_result217[95]^and_result217[96]^and_result217[97]^and_result217[98]^and_result217[99]^and_result217[100]^and_result217[101]^and_result217[102]^and_result217[103]^and_result217[104]^and_result217[105]^and_result217[106]^and_result217[107]^and_result217[108]^and_result217[109]^and_result217[110]^and_result217[111]^and_result217[112]^and_result217[113]^and_result217[114]^and_result217[115]^and_result217[116]^and_result217[117]^and_result217[118]^and_result217[119]^and_result217[120]^and_result217[121]^and_result217[122]^and_result217[123]^and_result217[124]^and_result217[125]^and_result217[126]^and_result217[127]^and_result217[128]^and_result217[129]^and_result217[130]^and_result217[131]^and_result217[132]^and_result217[133]^and_result217[134]^and_result217[135]^and_result217[136]^and_result217[137]^and_result217[138]^and_result217[139]^and_result217[140]^and_result217[141]^and_result217[142]^and_result217[143]^and_result217[144]^and_result217[145]^and_result217[146]^and_result217[147]^and_result217[148]^and_result217[149]^and_result217[150]^and_result217[151]^and_result217[152]^and_result217[153]^and_result217[154]^and_result217[155]^and_result217[156]^and_result217[157]^and_result217[158]^and_result217[159]^and_result217[160]^and_result217[161]^and_result217[162]^and_result217[163]^and_result217[164]^and_result217[165]^and_result217[166]^and_result217[167]^and_result217[168]^and_result217[169]^and_result217[170]^and_result217[171]^and_result217[172]^and_result217[173]^and_result217[174]^and_result217[175]^and_result217[176]^and_result217[177]^and_result217[178]^and_result217[179]^and_result217[180]^and_result217[181]^and_result217[182]^and_result217[183]^and_result217[184]^and_result217[185]^and_result217[186]^and_result217[187]^and_result217[188]^and_result217[189]^and_result217[190]^and_result217[191]^and_result217[192]^and_result217[193]^and_result217[194]^and_result217[195]^and_result217[196]^and_result217[197]^and_result217[198]^and_result217[199]^and_result217[200]^and_result217[201]^and_result217[202]^and_result217[203]^and_result217[204]^and_result217[205]^and_result217[206]^and_result217[207]^and_result217[208]^and_result217[209]^and_result217[210]^and_result217[211]^and_result217[212]^and_result217[213]^and_result217[214]^and_result217[215]^and_result217[216]^and_result217[217]^and_result217[218]^and_result217[219]^and_result217[220]^and_result217[221]^and_result217[222]^and_result217[223]^and_result217[224]^and_result217[225]^and_result217[226]^and_result217[227]^and_result217[228]^and_result217[229]^and_result217[230]^and_result217[231]^and_result217[232]^and_result217[233]^and_result217[234]^and_result217[235]^and_result217[236]^and_result217[237]^and_result217[238]^and_result217[239]^and_result217[240]^and_result217[241]^and_result217[242]^and_result217[243]^and_result217[244]^and_result217[245]^and_result217[246]^and_result217[247]^and_result217[248]^and_result217[249]^and_result217[250]^and_result217[251]^and_result217[252]^and_result217[253]^and_result217[254];
assign key[218]=and_result218[0]^and_result218[1]^and_result218[2]^and_result218[3]^and_result218[4]^and_result218[5]^and_result218[6]^and_result218[7]^and_result218[8]^and_result218[9]^and_result218[10]^and_result218[11]^and_result218[12]^and_result218[13]^and_result218[14]^and_result218[15]^and_result218[16]^and_result218[17]^and_result218[18]^and_result218[19]^and_result218[20]^and_result218[21]^and_result218[22]^and_result218[23]^and_result218[24]^and_result218[25]^and_result218[26]^and_result218[27]^and_result218[28]^and_result218[29]^and_result218[30]^and_result218[31]^and_result218[32]^and_result218[33]^and_result218[34]^and_result218[35]^and_result218[36]^and_result218[37]^and_result218[38]^and_result218[39]^and_result218[40]^and_result218[41]^and_result218[42]^and_result218[43]^and_result218[44]^and_result218[45]^and_result218[46]^and_result218[47]^and_result218[48]^and_result218[49]^and_result218[50]^and_result218[51]^and_result218[52]^and_result218[53]^and_result218[54]^and_result218[55]^and_result218[56]^and_result218[57]^and_result218[58]^and_result218[59]^and_result218[60]^and_result218[61]^and_result218[62]^and_result218[63]^and_result218[64]^and_result218[65]^and_result218[66]^and_result218[67]^and_result218[68]^and_result218[69]^and_result218[70]^and_result218[71]^and_result218[72]^and_result218[73]^and_result218[74]^and_result218[75]^and_result218[76]^and_result218[77]^and_result218[78]^and_result218[79]^and_result218[80]^and_result218[81]^and_result218[82]^and_result218[83]^and_result218[84]^and_result218[85]^and_result218[86]^and_result218[87]^and_result218[88]^and_result218[89]^and_result218[90]^and_result218[91]^and_result218[92]^and_result218[93]^and_result218[94]^and_result218[95]^and_result218[96]^and_result218[97]^and_result218[98]^and_result218[99]^and_result218[100]^and_result218[101]^and_result218[102]^and_result218[103]^and_result218[104]^and_result218[105]^and_result218[106]^and_result218[107]^and_result218[108]^and_result218[109]^and_result218[110]^and_result218[111]^and_result218[112]^and_result218[113]^and_result218[114]^and_result218[115]^and_result218[116]^and_result218[117]^and_result218[118]^and_result218[119]^and_result218[120]^and_result218[121]^and_result218[122]^and_result218[123]^and_result218[124]^and_result218[125]^and_result218[126]^and_result218[127]^and_result218[128]^and_result218[129]^and_result218[130]^and_result218[131]^and_result218[132]^and_result218[133]^and_result218[134]^and_result218[135]^and_result218[136]^and_result218[137]^and_result218[138]^and_result218[139]^and_result218[140]^and_result218[141]^and_result218[142]^and_result218[143]^and_result218[144]^and_result218[145]^and_result218[146]^and_result218[147]^and_result218[148]^and_result218[149]^and_result218[150]^and_result218[151]^and_result218[152]^and_result218[153]^and_result218[154]^and_result218[155]^and_result218[156]^and_result218[157]^and_result218[158]^and_result218[159]^and_result218[160]^and_result218[161]^and_result218[162]^and_result218[163]^and_result218[164]^and_result218[165]^and_result218[166]^and_result218[167]^and_result218[168]^and_result218[169]^and_result218[170]^and_result218[171]^and_result218[172]^and_result218[173]^and_result218[174]^and_result218[175]^and_result218[176]^and_result218[177]^and_result218[178]^and_result218[179]^and_result218[180]^and_result218[181]^and_result218[182]^and_result218[183]^and_result218[184]^and_result218[185]^and_result218[186]^and_result218[187]^and_result218[188]^and_result218[189]^and_result218[190]^and_result218[191]^and_result218[192]^and_result218[193]^and_result218[194]^and_result218[195]^and_result218[196]^and_result218[197]^and_result218[198]^and_result218[199]^and_result218[200]^and_result218[201]^and_result218[202]^and_result218[203]^and_result218[204]^and_result218[205]^and_result218[206]^and_result218[207]^and_result218[208]^and_result218[209]^and_result218[210]^and_result218[211]^and_result218[212]^and_result218[213]^and_result218[214]^and_result218[215]^and_result218[216]^and_result218[217]^and_result218[218]^and_result218[219]^and_result218[220]^and_result218[221]^and_result218[222]^and_result218[223]^and_result218[224]^and_result218[225]^and_result218[226]^and_result218[227]^and_result218[228]^and_result218[229]^and_result218[230]^and_result218[231]^and_result218[232]^and_result218[233]^and_result218[234]^and_result218[235]^and_result218[236]^and_result218[237]^and_result218[238]^and_result218[239]^and_result218[240]^and_result218[241]^and_result218[242]^and_result218[243]^and_result218[244]^and_result218[245]^and_result218[246]^and_result218[247]^and_result218[248]^and_result218[249]^and_result218[250]^and_result218[251]^and_result218[252]^and_result218[253]^and_result218[254];
assign key[219]=and_result219[0]^and_result219[1]^and_result219[2]^and_result219[3]^and_result219[4]^and_result219[5]^and_result219[6]^and_result219[7]^and_result219[8]^and_result219[9]^and_result219[10]^and_result219[11]^and_result219[12]^and_result219[13]^and_result219[14]^and_result219[15]^and_result219[16]^and_result219[17]^and_result219[18]^and_result219[19]^and_result219[20]^and_result219[21]^and_result219[22]^and_result219[23]^and_result219[24]^and_result219[25]^and_result219[26]^and_result219[27]^and_result219[28]^and_result219[29]^and_result219[30]^and_result219[31]^and_result219[32]^and_result219[33]^and_result219[34]^and_result219[35]^and_result219[36]^and_result219[37]^and_result219[38]^and_result219[39]^and_result219[40]^and_result219[41]^and_result219[42]^and_result219[43]^and_result219[44]^and_result219[45]^and_result219[46]^and_result219[47]^and_result219[48]^and_result219[49]^and_result219[50]^and_result219[51]^and_result219[52]^and_result219[53]^and_result219[54]^and_result219[55]^and_result219[56]^and_result219[57]^and_result219[58]^and_result219[59]^and_result219[60]^and_result219[61]^and_result219[62]^and_result219[63]^and_result219[64]^and_result219[65]^and_result219[66]^and_result219[67]^and_result219[68]^and_result219[69]^and_result219[70]^and_result219[71]^and_result219[72]^and_result219[73]^and_result219[74]^and_result219[75]^and_result219[76]^and_result219[77]^and_result219[78]^and_result219[79]^and_result219[80]^and_result219[81]^and_result219[82]^and_result219[83]^and_result219[84]^and_result219[85]^and_result219[86]^and_result219[87]^and_result219[88]^and_result219[89]^and_result219[90]^and_result219[91]^and_result219[92]^and_result219[93]^and_result219[94]^and_result219[95]^and_result219[96]^and_result219[97]^and_result219[98]^and_result219[99]^and_result219[100]^and_result219[101]^and_result219[102]^and_result219[103]^and_result219[104]^and_result219[105]^and_result219[106]^and_result219[107]^and_result219[108]^and_result219[109]^and_result219[110]^and_result219[111]^and_result219[112]^and_result219[113]^and_result219[114]^and_result219[115]^and_result219[116]^and_result219[117]^and_result219[118]^and_result219[119]^and_result219[120]^and_result219[121]^and_result219[122]^and_result219[123]^and_result219[124]^and_result219[125]^and_result219[126]^and_result219[127]^and_result219[128]^and_result219[129]^and_result219[130]^and_result219[131]^and_result219[132]^and_result219[133]^and_result219[134]^and_result219[135]^and_result219[136]^and_result219[137]^and_result219[138]^and_result219[139]^and_result219[140]^and_result219[141]^and_result219[142]^and_result219[143]^and_result219[144]^and_result219[145]^and_result219[146]^and_result219[147]^and_result219[148]^and_result219[149]^and_result219[150]^and_result219[151]^and_result219[152]^and_result219[153]^and_result219[154]^and_result219[155]^and_result219[156]^and_result219[157]^and_result219[158]^and_result219[159]^and_result219[160]^and_result219[161]^and_result219[162]^and_result219[163]^and_result219[164]^and_result219[165]^and_result219[166]^and_result219[167]^and_result219[168]^and_result219[169]^and_result219[170]^and_result219[171]^and_result219[172]^and_result219[173]^and_result219[174]^and_result219[175]^and_result219[176]^and_result219[177]^and_result219[178]^and_result219[179]^and_result219[180]^and_result219[181]^and_result219[182]^and_result219[183]^and_result219[184]^and_result219[185]^and_result219[186]^and_result219[187]^and_result219[188]^and_result219[189]^and_result219[190]^and_result219[191]^and_result219[192]^and_result219[193]^and_result219[194]^and_result219[195]^and_result219[196]^and_result219[197]^and_result219[198]^and_result219[199]^and_result219[200]^and_result219[201]^and_result219[202]^and_result219[203]^and_result219[204]^and_result219[205]^and_result219[206]^and_result219[207]^and_result219[208]^and_result219[209]^and_result219[210]^and_result219[211]^and_result219[212]^and_result219[213]^and_result219[214]^and_result219[215]^and_result219[216]^and_result219[217]^and_result219[218]^and_result219[219]^and_result219[220]^and_result219[221]^and_result219[222]^and_result219[223]^and_result219[224]^and_result219[225]^and_result219[226]^and_result219[227]^and_result219[228]^and_result219[229]^and_result219[230]^and_result219[231]^and_result219[232]^and_result219[233]^and_result219[234]^and_result219[235]^and_result219[236]^and_result219[237]^and_result219[238]^and_result219[239]^and_result219[240]^and_result219[241]^and_result219[242]^and_result219[243]^and_result219[244]^and_result219[245]^and_result219[246]^and_result219[247]^and_result219[248]^and_result219[249]^and_result219[250]^and_result219[251]^and_result219[252]^and_result219[253]^and_result219[254];
assign key[220]=and_result220[0]^and_result220[1]^and_result220[2]^and_result220[3]^and_result220[4]^and_result220[5]^and_result220[6]^and_result220[7]^and_result220[8]^and_result220[9]^and_result220[10]^and_result220[11]^and_result220[12]^and_result220[13]^and_result220[14]^and_result220[15]^and_result220[16]^and_result220[17]^and_result220[18]^and_result220[19]^and_result220[20]^and_result220[21]^and_result220[22]^and_result220[23]^and_result220[24]^and_result220[25]^and_result220[26]^and_result220[27]^and_result220[28]^and_result220[29]^and_result220[30]^and_result220[31]^and_result220[32]^and_result220[33]^and_result220[34]^and_result220[35]^and_result220[36]^and_result220[37]^and_result220[38]^and_result220[39]^and_result220[40]^and_result220[41]^and_result220[42]^and_result220[43]^and_result220[44]^and_result220[45]^and_result220[46]^and_result220[47]^and_result220[48]^and_result220[49]^and_result220[50]^and_result220[51]^and_result220[52]^and_result220[53]^and_result220[54]^and_result220[55]^and_result220[56]^and_result220[57]^and_result220[58]^and_result220[59]^and_result220[60]^and_result220[61]^and_result220[62]^and_result220[63]^and_result220[64]^and_result220[65]^and_result220[66]^and_result220[67]^and_result220[68]^and_result220[69]^and_result220[70]^and_result220[71]^and_result220[72]^and_result220[73]^and_result220[74]^and_result220[75]^and_result220[76]^and_result220[77]^and_result220[78]^and_result220[79]^and_result220[80]^and_result220[81]^and_result220[82]^and_result220[83]^and_result220[84]^and_result220[85]^and_result220[86]^and_result220[87]^and_result220[88]^and_result220[89]^and_result220[90]^and_result220[91]^and_result220[92]^and_result220[93]^and_result220[94]^and_result220[95]^and_result220[96]^and_result220[97]^and_result220[98]^and_result220[99]^and_result220[100]^and_result220[101]^and_result220[102]^and_result220[103]^and_result220[104]^and_result220[105]^and_result220[106]^and_result220[107]^and_result220[108]^and_result220[109]^and_result220[110]^and_result220[111]^and_result220[112]^and_result220[113]^and_result220[114]^and_result220[115]^and_result220[116]^and_result220[117]^and_result220[118]^and_result220[119]^and_result220[120]^and_result220[121]^and_result220[122]^and_result220[123]^and_result220[124]^and_result220[125]^and_result220[126]^and_result220[127]^and_result220[128]^and_result220[129]^and_result220[130]^and_result220[131]^and_result220[132]^and_result220[133]^and_result220[134]^and_result220[135]^and_result220[136]^and_result220[137]^and_result220[138]^and_result220[139]^and_result220[140]^and_result220[141]^and_result220[142]^and_result220[143]^and_result220[144]^and_result220[145]^and_result220[146]^and_result220[147]^and_result220[148]^and_result220[149]^and_result220[150]^and_result220[151]^and_result220[152]^and_result220[153]^and_result220[154]^and_result220[155]^and_result220[156]^and_result220[157]^and_result220[158]^and_result220[159]^and_result220[160]^and_result220[161]^and_result220[162]^and_result220[163]^and_result220[164]^and_result220[165]^and_result220[166]^and_result220[167]^and_result220[168]^and_result220[169]^and_result220[170]^and_result220[171]^and_result220[172]^and_result220[173]^and_result220[174]^and_result220[175]^and_result220[176]^and_result220[177]^and_result220[178]^and_result220[179]^and_result220[180]^and_result220[181]^and_result220[182]^and_result220[183]^and_result220[184]^and_result220[185]^and_result220[186]^and_result220[187]^and_result220[188]^and_result220[189]^and_result220[190]^and_result220[191]^and_result220[192]^and_result220[193]^and_result220[194]^and_result220[195]^and_result220[196]^and_result220[197]^and_result220[198]^and_result220[199]^and_result220[200]^and_result220[201]^and_result220[202]^and_result220[203]^and_result220[204]^and_result220[205]^and_result220[206]^and_result220[207]^and_result220[208]^and_result220[209]^and_result220[210]^and_result220[211]^and_result220[212]^and_result220[213]^and_result220[214]^and_result220[215]^and_result220[216]^and_result220[217]^and_result220[218]^and_result220[219]^and_result220[220]^and_result220[221]^and_result220[222]^and_result220[223]^and_result220[224]^and_result220[225]^and_result220[226]^and_result220[227]^and_result220[228]^and_result220[229]^and_result220[230]^and_result220[231]^and_result220[232]^and_result220[233]^and_result220[234]^and_result220[235]^and_result220[236]^and_result220[237]^and_result220[238]^and_result220[239]^and_result220[240]^and_result220[241]^and_result220[242]^and_result220[243]^and_result220[244]^and_result220[245]^and_result220[246]^and_result220[247]^and_result220[248]^and_result220[249]^and_result220[250]^and_result220[251]^and_result220[252]^and_result220[253]^and_result220[254];
assign key[221]=and_result221[0]^and_result221[1]^and_result221[2]^and_result221[3]^and_result221[4]^and_result221[5]^and_result221[6]^and_result221[7]^and_result221[8]^and_result221[9]^and_result221[10]^and_result221[11]^and_result221[12]^and_result221[13]^and_result221[14]^and_result221[15]^and_result221[16]^and_result221[17]^and_result221[18]^and_result221[19]^and_result221[20]^and_result221[21]^and_result221[22]^and_result221[23]^and_result221[24]^and_result221[25]^and_result221[26]^and_result221[27]^and_result221[28]^and_result221[29]^and_result221[30]^and_result221[31]^and_result221[32]^and_result221[33]^and_result221[34]^and_result221[35]^and_result221[36]^and_result221[37]^and_result221[38]^and_result221[39]^and_result221[40]^and_result221[41]^and_result221[42]^and_result221[43]^and_result221[44]^and_result221[45]^and_result221[46]^and_result221[47]^and_result221[48]^and_result221[49]^and_result221[50]^and_result221[51]^and_result221[52]^and_result221[53]^and_result221[54]^and_result221[55]^and_result221[56]^and_result221[57]^and_result221[58]^and_result221[59]^and_result221[60]^and_result221[61]^and_result221[62]^and_result221[63]^and_result221[64]^and_result221[65]^and_result221[66]^and_result221[67]^and_result221[68]^and_result221[69]^and_result221[70]^and_result221[71]^and_result221[72]^and_result221[73]^and_result221[74]^and_result221[75]^and_result221[76]^and_result221[77]^and_result221[78]^and_result221[79]^and_result221[80]^and_result221[81]^and_result221[82]^and_result221[83]^and_result221[84]^and_result221[85]^and_result221[86]^and_result221[87]^and_result221[88]^and_result221[89]^and_result221[90]^and_result221[91]^and_result221[92]^and_result221[93]^and_result221[94]^and_result221[95]^and_result221[96]^and_result221[97]^and_result221[98]^and_result221[99]^and_result221[100]^and_result221[101]^and_result221[102]^and_result221[103]^and_result221[104]^and_result221[105]^and_result221[106]^and_result221[107]^and_result221[108]^and_result221[109]^and_result221[110]^and_result221[111]^and_result221[112]^and_result221[113]^and_result221[114]^and_result221[115]^and_result221[116]^and_result221[117]^and_result221[118]^and_result221[119]^and_result221[120]^and_result221[121]^and_result221[122]^and_result221[123]^and_result221[124]^and_result221[125]^and_result221[126]^and_result221[127]^and_result221[128]^and_result221[129]^and_result221[130]^and_result221[131]^and_result221[132]^and_result221[133]^and_result221[134]^and_result221[135]^and_result221[136]^and_result221[137]^and_result221[138]^and_result221[139]^and_result221[140]^and_result221[141]^and_result221[142]^and_result221[143]^and_result221[144]^and_result221[145]^and_result221[146]^and_result221[147]^and_result221[148]^and_result221[149]^and_result221[150]^and_result221[151]^and_result221[152]^and_result221[153]^and_result221[154]^and_result221[155]^and_result221[156]^and_result221[157]^and_result221[158]^and_result221[159]^and_result221[160]^and_result221[161]^and_result221[162]^and_result221[163]^and_result221[164]^and_result221[165]^and_result221[166]^and_result221[167]^and_result221[168]^and_result221[169]^and_result221[170]^and_result221[171]^and_result221[172]^and_result221[173]^and_result221[174]^and_result221[175]^and_result221[176]^and_result221[177]^and_result221[178]^and_result221[179]^and_result221[180]^and_result221[181]^and_result221[182]^and_result221[183]^and_result221[184]^and_result221[185]^and_result221[186]^and_result221[187]^and_result221[188]^and_result221[189]^and_result221[190]^and_result221[191]^and_result221[192]^and_result221[193]^and_result221[194]^and_result221[195]^and_result221[196]^and_result221[197]^and_result221[198]^and_result221[199]^and_result221[200]^and_result221[201]^and_result221[202]^and_result221[203]^and_result221[204]^and_result221[205]^and_result221[206]^and_result221[207]^and_result221[208]^and_result221[209]^and_result221[210]^and_result221[211]^and_result221[212]^and_result221[213]^and_result221[214]^and_result221[215]^and_result221[216]^and_result221[217]^and_result221[218]^and_result221[219]^and_result221[220]^and_result221[221]^and_result221[222]^and_result221[223]^and_result221[224]^and_result221[225]^and_result221[226]^and_result221[227]^and_result221[228]^and_result221[229]^and_result221[230]^and_result221[231]^and_result221[232]^and_result221[233]^and_result221[234]^and_result221[235]^and_result221[236]^and_result221[237]^and_result221[238]^and_result221[239]^and_result221[240]^and_result221[241]^and_result221[242]^and_result221[243]^and_result221[244]^and_result221[245]^and_result221[246]^and_result221[247]^and_result221[248]^and_result221[249]^and_result221[250]^and_result221[251]^and_result221[252]^and_result221[253]^and_result221[254];
assign key[222]=and_result222[0]^and_result222[1]^and_result222[2]^and_result222[3]^and_result222[4]^and_result222[5]^and_result222[6]^and_result222[7]^and_result222[8]^and_result222[9]^and_result222[10]^and_result222[11]^and_result222[12]^and_result222[13]^and_result222[14]^and_result222[15]^and_result222[16]^and_result222[17]^and_result222[18]^and_result222[19]^and_result222[20]^and_result222[21]^and_result222[22]^and_result222[23]^and_result222[24]^and_result222[25]^and_result222[26]^and_result222[27]^and_result222[28]^and_result222[29]^and_result222[30]^and_result222[31]^and_result222[32]^and_result222[33]^and_result222[34]^and_result222[35]^and_result222[36]^and_result222[37]^and_result222[38]^and_result222[39]^and_result222[40]^and_result222[41]^and_result222[42]^and_result222[43]^and_result222[44]^and_result222[45]^and_result222[46]^and_result222[47]^and_result222[48]^and_result222[49]^and_result222[50]^and_result222[51]^and_result222[52]^and_result222[53]^and_result222[54]^and_result222[55]^and_result222[56]^and_result222[57]^and_result222[58]^and_result222[59]^and_result222[60]^and_result222[61]^and_result222[62]^and_result222[63]^and_result222[64]^and_result222[65]^and_result222[66]^and_result222[67]^and_result222[68]^and_result222[69]^and_result222[70]^and_result222[71]^and_result222[72]^and_result222[73]^and_result222[74]^and_result222[75]^and_result222[76]^and_result222[77]^and_result222[78]^and_result222[79]^and_result222[80]^and_result222[81]^and_result222[82]^and_result222[83]^and_result222[84]^and_result222[85]^and_result222[86]^and_result222[87]^and_result222[88]^and_result222[89]^and_result222[90]^and_result222[91]^and_result222[92]^and_result222[93]^and_result222[94]^and_result222[95]^and_result222[96]^and_result222[97]^and_result222[98]^and_result222[99]^and_result222[100]^and_result222[101]^and_result222[102]^and_result222[103]^and_result222[104]^and_result222[105]^and_result222[106]^and_result222[107]^and_result222[108]^and_result222[109]^and_result222[110]^and_result222[111]^and_result222[112]^and_result222[113]^and_result222[114]^and_result222[115]^and_result222[116]^and_result222[117]^and_result222[118]^and_result222[119]^and_result222[120]^and_result222[121]^and_result222[122]^and_result222[123]^and_result222[124]^and_result222[125]^and_result222[126]^and_result222[127]^and_result222[128]^and_result222[129]^and_result222[130]^and_result222[131]^and_result222[132]^and_result222[133]^and_result222[134]^and_result222[135]^and_result222[136]^and_result222[137]^and_result222[138]^and_result222[139]^and_result222[140]^and_result222[141]^and_result222[142]^and_result222[143]^and_result222[144]^and_result222[145]^and_result222[146]^and_result222[147]^and_result222[148]^and_result222[149]^and_result222[150]^and_result222[151]^and_result222[152]^and_result222[153]^and_result222[154]^and_result222[155]^and_result222[156]^and_result222[157]^and_result222[158]^and_result222[159]^and_result222[160]^and_result222[161]^and_result222[162]^and_result222[163]^and_result222[164]^and_result222[165]^and_result222[166]^and_result222[167]^and_result222[168]^and_result222[169]^and_result222[170]^and_result222[171]^and_result222[172]^and_result222[173]^and_result222[174]^and_result222[175]^and_result222[176]^and_result222[177]^and_result222[178]^and_result222[179]^and_result222[180]^and_result222[181]^and_result222[182]^and_result222[183]^and_result222[184]^and_result222[185]^and_result222[186]^and_result222[187]^and_result222[188]^and_result222[189]^and_result222[190]^and_result222[191]^and_result222[192]^and_result222[193]^and_result222[194]^and_result222[195]^and_result222[196]^and_result222[197]^and_result222[198]^and_result222[199]^and_result222[200]^and_result222[201]^and_result222[202]^and_result222[203]^and_result222[204]^and_result222[205]^and_result222[206]^and_result222[207]^and_result222[208]^and_result222[209]^and_result222[210]^and_result222[211]^and_result222[212]^and_result222[213]^and_result222[214]^and_result222[215]^and_result222[216]^and_result222[217]^and_result222[218]^and_result222[219]^and_result222[220]^and_result222[221]^and_result222[222]^and_result222[223]^and_result222[224]^and_result222[225]^and_result222[226]^and_result222[227]^and_result222[228]^and_result222[229]^and_result222[230]^and_result222[231]^and_result222[232]^and_result222[233]^and_result222[234]^and_result222[235]^and_result222[236]^and_result222[237]^and_result222[238]^and_result222[239]^and_result222[240]^and_result222[241]^and_result222[242]^and_result222[243]^and_result222[244]^and_result222[245]^and_result222[246]^and_result222[247]^and_result222[248]^and_result222[249]^and_result222[250]^and_result222[251]^and_result222[252]^and_result222[253]^and_result222[254];
assign key[223]=and_result223[0]^and_result223[1]^and_result223[2]^and_result223[3]^and_result223[4]^and_result223[5]^and_result223[6]^and_result223[7]^and_result223[8]^and_result223[9]^and_result223[10]^and_result223[11]^and_result223[12]^and_result223[13]^and_result223[14]^and_result223[15]^and_result223[16]^and_result223[17]^and_result223[18]^and_result223[19]^and_result223[20]^and_result223[21]^and_result223[22]^and_result223[23]^and_result223[24]^and_result223[25]^and_result223[26]^and_result223[27]^and_result223[28]^and_result223[29]^and_result223[30]^and_result223[31]^and_result223[32]^and_result223[33]^and_result223[34]^and_result223[35]^and_result223[36]^and_result223[37]^and_result223[38]^and_result223[39]^and_result223[40]^and_result223[41]^and_result223[42]^and_result223[43]^and_result223[44]^and_result223[45]^and_result223[46]^and_result223[47]^and_result223[48]^and_result223[49]^and_result223[50]^and_result223[51]^and_result223[52]^and_result223[53]^and_result223[54]^and_result223[55]^and_result223[56]^and_result223[57]^and_result223[58]^and_result223[59]^and_result223[60]^and_result223[61]^and_result223[62]^and_result223[63]^and_result223[64]^and_result223[65]^and_result223[66]^and_result223[67]^and_result223[68]^and_result223[69]^and_result223[70]^and_result223[71]^and_result223[72]^and_result223[73]^and_result223[74]^and_result223[75]^and_result223[76]^and_result223[77]^and_result223[78]^and_result223[79]^and_result223[80]^and_result223[81]^and_result223[82]^and_result223[83]^and_result223[84]^and_result223[85]^and_result223[86]^and_result223[87]^and_result223[88]^and_result223[89]^and_result223[90]^and_result223[91]^and_result223[92]^and_result223[93]^and_result223[94]^and_result223[95]^and_result223[96]^and_result223[97]^and_result223[98]^and_result223[99]^and_result223[100]^and_result223[101]^and_result223[102]^and_result223[103]^and_result223[104]^and_result223[105]^and_result223[106]^and_result223[107]^and_result223[108]^and_result223[109]^and_result223[110]^and_result223[111]^and_result223[112]^and_result223[113]^and_result223[114]^and_result223[115]^and_result223[116]^and_result223[117]^and_result223[118]^and_result223[119]^and_result223[120]^and_result223[121]^and_result223[122]^and_result223[123]^and_result223[124]^and_result223[125]^and_result223[126]^and_result223[127]^and_result223[128]^and_result223[129]^and_result223[130]^and_result223[131]^and_result223[132]^and_result223[133]^and_result223[134]^and_result223[135]^and_result223[136]^and_result223[137]^and_result223[138]^and_result223[139]^and_result223[140]^and_result223[141]^and_result223[142]^and_result223[143]^and_result223[144]^and_result223[145]^and_result223[146]^and_result223[147]^and_result223[148]^and_result223[149]^and_result223[150]^and_result223[151]^and_result223[152]^and_result223[153]^and_result223[154]^and_result223[155]^and_result223[156]^and_result223[157]^and_result223[158]^and_result223[159]^and_result223[160]^and_result223[161]^and_result223[162]^and_result223[163]^and_result223[164]^and_result223[165]^and_result223[166]^and_result223[167]^and_result223[168]^and_result223[169]^and_result223[170]^and_result223[171]^and_result223[172]^and_result223[173]^and_result223[174]^and_result223[175]^and_result223[176]^and_result223[177]^and_result223[178]^and_result223[179]^and_result223[180]^and_result223[181]^and_result223[182]^and_result223[183]^and_result223[184]^and_result223[185]^and_result223[186]^and_result223[187]^and_result223[188]^and_result223[189]^and_result223[190]^and_result223[191]^and_result223[192]^and_result223[193]^and_result223[194]^and_result223[195]^and_result223[196]^and_result223[197]^and_result223[198]^and_result223[199]^and_result223[200]^and_result223[201]^and_result223[202]^and_result223[203]^and_result223[204]^and_result223[205]^and_result223[206]^and_result223[207]^and_result223[208]^and_result223[209]^and_result223[210]^and_result223[211]^and_result223[212]^and_result223[213]^and_result223[214]^and_result223[215]^and_result223[216]^and_result223[217]^and_result223[218]^and_result223[219]^and_result223[220]^and_result223[221]^and_result223[222]^and_result223[223]^and_result223[224]^and_result223[225]^and_result223[226]^and_result223[227]^and_result223[228]^and_result223[229]^and_result223[230]^and_result223[231]^and_result223[232]^and_result223[233]^and_result223[234]^and_result223[235]^and_result223[236]^and_result223[237]^and_result223[238]^and_result223[239]^and_result223[240]^and_result223[241]^and_result223[242]^and_result223[243]^and_result223[244]^and_result223[245]^and_result223[246]^and_result223[247]^and_result223[248]^and_result223[249]^and_result223[250]^and_result223[251]^and_result223[252]^and_result223[253]^and_result223[254];
assign key[224]=and_result224[0]^and_result224[1]^and_result224[2]^and_result224[3]^and_result224[4]^and_result224[5]^and_result224[6]^and_result224[7]^and_result224[8]^and_result224[9]^and_result224[10]^and_result224[11]^and_result224[12]^and_result224[13]^and_result224[14]^and_result224[15]^and_result224[16]^and_result224[17]^and_result224[18]^and_result224[19]^and_result224[20]^and_result224[21]^and_result224[22]^and_result224[23]^and_result224[24]^and_result224[25]^and_result224[26]^and_result224[27]^and_result224[28]^and_result224[29]^and_result224[30]^and_result224[31]^and_result224[32]^and_result224[33]^and_result224[34]^and_result224[35]^and_result224[36]^and_result224[37]^and_result224[38]^and_result224[39]^and_result224[40]^and_result224[41]^and_result224[42]^and_result224[43]^and_result224[44]^and_result224[45]^and_result224[46]^and_result224[47]^and_result224[48]^and_result224[49]^and_result224[50]^and_result224[51]^and_result224[52]^and_result224[53]^and_result224[54]^and_result224[55]^and_result224[56]^and_result224[57]^and_result224[58]^and_result224[59]^and_result224[60]^and_result224[61]^and_result224[62]^and_result224[63]^and_result224[64]^and_result224[65]^and_result224[66]^and_result224[67]^and_result224[68]^and_result224[69]^and_result224[70]^and_result224[71]^and_result224[72]^and_result224[73]^and_result224[74]^and_result224[75]^and_result224[76]^and_result224[77]^and_result224[78]^and_result224[79]^and_result224[80]^and_result224[81]^and_result224[82]^and_result224[83]^and_result224[84]^and_result224[85]^and_result224[86]^and_result224[87]^and_result224[88]^and_result224[89]^and_result224[90]^and_result224[91]^and_result224[92]^and_result224[93]^and_result224[94]^and_result224[95]^and_result224[96]^and_result224[97]^and_result224[98]^and_result224[99]^and_result224[100]^and_result224[101]^and_result224[102]^and_result224[103]^and_result224[104]^and_result224[105]^and_result224[106]^and_result224[107]^and_result224[108]^and_result224[109]^and_result224[110]^and_result224[111]^and_result224[112]^and_result224[113]^and_result224[114]^and_result224[115]^and_result224[116]^and_result224[117]^and_result224[118]^and_result224[119]^and_result224[120]^and_result224[121]^and_result224[122]^and_result224[123]^and_result224[124]^and_result224[125]^and_result224[126]^and_result224[127]^and_result224[128]^and_result224[129]^and_result224[130]^and_result224[131]^and_result224[132]^and_result224[133]^and_result224[134]^and_result224[135]^and_result224[136]^and_result224[137]^and_result224[138]^and_result224[139]^and_result224[140]^and_result224[141]^and_result224[142]^and_result224[143]^and_result224[144]^and_result224[145]^and_result224[146]^and_result224[147]^and_result224[148]^and_result224[149]^and_result224[150]^and_result224[151]^and_result224[152]^and_result224[153]^and_result224[154]^and_result224[155]^and_result224[156]^and_result224[157]^and_result224[158]^and_result224[159]^and_result224[160]^and_result224[161]^and_result224[162]^and_result224[163]^and_result224[164]^and_result224[165]^and_result224[166]^and_result224[167]^and_result224[168]^and_result224[169]^and_result224[170]^and_result224[171]^and_result224[172]^and_result224[173]^and_result224[174]^and_result224[175]^and_result224[176]^and_result224[177]^and_result224[178]^and_result224[179]^and_result224[180]^and_result224[181]^and_result224[182]^and_result224[183]^and_result224[184]^and_result224[185]^and_result224[186]^and_result224[187]^and_result224[188]^and_result224[189]^and_result224[190]^and_result224[191]^and_result224[192]^and_result224[193]^and_result224[194]^and_result224[195]^and_result224[196]^and_result224[197]^and_result224[198]^and_result224[199]^and_result224[200]^and_result224[201]^and_result224[202]^and_result224[203]^and_result224[204]^and_result224[205]^and_result224[206]^and_result224[207]^and_result224[208]^and_result224[209]^and_result224[210]^and_result224[211]^and_result224[212]^and_result224[213]^and_result224[214]^and_result224[215]^and_result224[216]^and_result224[217]^and_result224[218]^and_result224[219]^and_result224[220]^and_result224[221]^and_result224[222]^and_result224[223]^and_result224[224]^and_result224[225]^and_result224[226]^and_result224[227]^and_result224[228]^and_result224[229]^and_result224[230]^and_result224[231]^and_result224[232]^and_result224[233]^and_result224[234]^and_result224[235]^and_result224[236]^and_result224[237]^and_result224[238]^and_result224[239]^and_result224[240]^and_result224[241]^and_result224[242]^and_result224[243]^and_result224[244]^and_result224[245]^and_result224[246]^and_result224[247]^and_result224[248]^and_result224[249]^and_result224[250]^and_result224[251]^and_result224[252]^and_result224[253]^and_result224[254];
assign key[225]=and_result225[0]^and_result225[1]^and_result225[2]^and_result225[3]^and_result225[4]^and_result225[5]^and_result225[6]^and_result225[7]^and_result225[8]^and_result225[9]^and_result225[10]^and_result225[11]^and_result225[12]^and_result225[13]^and_result225[14]^and_result225[15]^and_result225[16]^and_result225[17]^and_result225[18]^and_result225[19]^and_result225[20]^and_result225[21]^and_result225[22]^and_result225[23]^and_result225[24]^and_result225[25]^and_result225[26]^and_result225[27]^and_result225[28]^and_result225[29]^and_result225[30]^and_result225[31]^and_result225[32]^and_result225[33]^and_result225[34]^and_result225[35]^and_result225[36]^and_result225[37]^and_result225[38]^and_result225[39]^and_result225[40]^and_result225[41]^and_result225[42]^and_result225[43]^and_result225[44]^and_result225[45]^and_result225[46]^and_result225[47]^and_result225[48]^and_result225[49]^and_result225[50]^and_result225[51]^and_result225[52]^and_result225[53]^and_result225[54]^and_result225[55]^and_result225[56]^and_result225[57]^and_result225[58]^and_result225[59]^and_result225[60]^and_result225[61]^and_result225[62]^and_result225[63]^and_result225[64]^and_result225[65]^and_result225[66]^and_result225[67]^and_result225[68]^and_result225[69]^and_result225[70]^and_result225[71]^and_result225[72]^and_result225[73]^and_result225[74]^and_result225[75]^and_result225[76]^and_result225[77]^and_result225[78]^and_result225[79]^and_result225[80]^and_result225[81]^and_result225[82]^and_result225[83]^and_result225[84]^and_result225[85]^and_result225[86]^and_result225[87]^and_result225[88]^and_result225[89]^and_result225[90]^and_result225[91]^and_result225[92]^and_result225[93]^and_result225[94]^and_result225[95]^and_result225[96]^and_result225[97]^and_result225[98]^and_result225[99]^and_result225[100]^and_result225[101]^and_result225[102]^and_result225[103]^and_result225[104]^and_result225[105]^and_result225[106]^and_result225[107]^and_result225[108]^and_result225[109]^and_result225[110]^and_result225[111]^and_result225[112]^and_result225[113]^and_result225[114]^and_result225[115]^and_result225[116]^and_result225[117]^and_result225[118]^and_result225[119]^and_result225[120]^and_result225[121]^and_result225[122]^and_result225[123]^and_result225[124]^and_result225[125]^and_result225[126]^and_result225[127]^and_result225[128]^and_result225[129]^and_result225[130]^and_result225[131]^and_result225[132]^and_result225[133]^and_result225[134]^and_result225[135]^and_result225[136]^and_result225[137]^and_result225[138]^and_result225[139]^and_result225[140]^and_result225[141]^and_result225[142]^and_result225[143]^and_result225[144]^and_result225[145]^and_result225[146]^and_result225[147]^and_result225[148]^and_result225[149]^and_result225[150]^and_result225[151]^and_result225[152]^and_result225[153]^and_result225[154]^and_result225[155]^and_result225[156]^and_result225[157]^and_result225[158]^and_result225[159]^and_result225[160]^and_result225[161]^and_result225[162]^and_result225[163]^and_result225[164]^and_result225[165]^and_result225[166]^and_result225[167]^and_result225[168]^and_result225[169]^and_result225[170]^and_result225[171]^and_result225[172]^and_result225[173]^and_result225[174]^and_result225[175]^and_result225[176]^and_result225[177]^and_result225[178]^and_result225[179]^and_result225[180]^and_result225[181]^and_result225[182]^and_result225[183]^and_result225[184]^and_result225[185]^and_result225[186]^and_result225[187]^and_result225[188]^and_result225[189]^and_result225[190]^and_result225[191]^and_result225[192]^and_result225[193]^and_result225[194]^and_result225[195]^and_result225[196]^and_result225[197]^and_result225[198]^and_result225[199]^and_result225[200]^and_result225[201]^and_result225[202]^and_result225[203]^and_result225[204]^and_result225[205]^and_result225[206]^and_result225[207]^and_result225[208]^and_result225[209]^and_result225[210]^and_result225[211]^and_result225[212]^and_result225[213]^and_result225[214]^and_result225[215]^and_result225[216]^and_result225[217]^and_result225[218]^and_result225[219]^and_result225[220]^and_result225[221]^and_result225[222]^and_result225[223]^and_result225[224]^and_result225[225]^and_result225[226]^and_result225[227]^and_result225[228]^and_result225[229]^and_result225[230]^and_result225[231]^and_result225[232]^and_result225[233]^and_result225[234]^and_result225[235]^and_result225[236]^and_result225[237]^and_result225[238]^and_result225[239]^and_result225[240]^and_result225[241]^and_result225[242]^and_result225[243]^and_result225[244]^and_result225[245]^and_result225[246]^and_result225[247]^and_result225[248]^and_result225[249]^and_result225[250]^and_result225[251]^and_result225[252]^and_result225[253]^and_result225[254];
assign key[226]=and_result226[0]^and_result226[1]^and_result226[2]^and_result226[3]^and_result226[4]^and_result226[5]^and_result226[6]^and_result226[7]^and_result226[8]^and_result226[9]^and_result226[10]^and_result226[11]^and_result226[12]^and_result226[13]^and_result226[14]^and_result226[15]^and_result226[16]^and_result226[17]^and_result226[18]^and_result226[19]^and_result226[20]^and_result226[21]^and_result226[22]^and_result226[23]^and_result226[24]^and_result226[25]^and_result226[26]^and_result226[27]^and_result226[28]^and_result226[29]^and_result226[30]^and_result226[31]^and_result226[32]^and_result226[33]^and_result226[34]^and_result226[35]^and_result226[36]^and_result226[37]^and_result226[38]^and_result226[39]^and_result226[40]^and_result226[41]^and_result226[42]^and_result226[43]^and_result226[44]^and_result226[45]^and_result226[46]^and_result226[47]^and_result226[48]^and_result226[49]^and_result226[50]^and_result226[51]^and_result226[52]^and_result226[53]^and_result226[54]^and_result226[55]^and_result226[56]^and_result226[57]^and_result226[58]^and_result226[59]^and_result226[60]^and_result226[61]^and_result226[62]^and_result226[63]^and_result226[64]^and_result226[65]^and_result226[66]^and_result226[67]^and_result226[68]^and_result226[69]^and_result226[70]^and_result226[71]^and_result226[72]^and_result226[73]^and_result226[74]^and_result226[75]^and_result226[76]^and_result226[77]^and_result226[78]^and_result226[79]^and_result226[80]^and_result226[81]^and_result226[82]^and_result226[83]^and_result226[84]^and_result226[85]^and_result226[86]^and_result226[87]^and_result226[88]^and_result226[89]^and_result226[90]^and_result226[91]^and_result226[92]^and_result226[93]^and_result226[94]^and_result226[95]^and_result226[96]^and_result226[97]^and_result226[98]^and_result226[99]^and_result226[100]^and_result226[101]^and_result226[102]^and_result226[103]^and_result226[104]^and_result226[105]^and_result226[106]^and_result226[107]^and_result226[108]^and_result226[109]^and_result226[110]^and_result226[111]^and_result226[112]^and_result226[113]^and_result226[114]^and_result226[115]^and_result226[116]^and_result226[117]^and_result226[118]^and_result226[119]^and_result226[120]^and_result226[121]^and_result226[122]^and_result226[123]^and_result226[124]^and_result226[125]^and_result226[126]^and_result226[127]^and_result226[128]^and_result226[129]^and_result226[130]^and_result226[131]^and_result226[132]^and_result226[133]^and_result226[134]^and_result226[135]^and_result226[136]^and_result226[137]^and_result226[138]^and_result226[139]^and_result226[140]^and_result226[141]^and_result226[142]^and_result226[143]^and_result226[144]^and_result226[145]^and_result226[146]^and_result226[147]^and_result226[148]^and_result226[149]^and_result226[150]^and_result226[151]^and_result226[152]^and_result226[153]^and_result226[154]^and_result226[155]^and_result226[156]^and_result226[157]^and_result226[158]^and_result226[159]^and_result226[160]^and_result226[161]^and_result226[162]^and_result226[163]^and_result226[164]^and_result226[165]^and_result226[166]^and_result226[167]^and_result226[168]^and_result226[169]^and_result226[170]^and_result226[171]^and_result226[172]^and_result226[173]^and_result226[174]^and_result226[175]^and_result226[176]^and_result226[177]^and_result226[178]^and_result226[179]^and_result226[180]^and_result226[181]^and_result226[182]^and_result226[183]^and_result226[184]^and_result226[185]^and_result226[186]^and_result226[187]^and_result226[188]^and_result226[189]^and_result226[190]^and_result226[191]^and_result226[192]^and_result226[193]^and_result226[194]^and_result226[195]^and_result226[196]^and_result226[197]^and_result226[198]^and_result226[199]^and_result226[200]^and_result226[201]^and_result226[202]^and_result226[203]^and_result226[204]^and_result226[205]^and_result226[206]^and_result226[207]^and_result226[208]^and_result226[209]^and_result226[210]^and_result226[211]^and_result226[212]^and_result226[213]^and_result226[214]^and_result226[215]^and_result226[216]^and_result226[217]^and_result226[218]^and_result226[219]^and_result226[220]^and_result226[221]^and_result226[222]^and_result226[223]^and_result226[224]^and_result226[225]^and_result226[226]^and_result226[227]^and_result226[228]^and_result226[229]^and_result226[230]^and_result226[231]^and_result226[232]^and_result226[233]^and_result226[234]^and_result226[235]^and_result226[236]^and_result226[237]^and_result226[238]^and_result226[239]^and_result226[240]^and_result226[241]^and_result226[242]^and_result226[243]^and_result226[244]^and_result226[245]^and_result226[246]^and_result226[247]^and_result226[248]^and_result226[249]^and_result226[250]^and_result226[251]^and_result226[252]^and_result226[253]^and_result226[254];
assign key[227]=and_result227[0]^and_result227[1]^and_result227[2]^and_result227[3]^and_result227[4]^and_result227[5]^and_result227[6]^and_result227[7]^and_result227[8]^and_result227[9]^and_result227[10]^and_result227[11]^and_result227[12]^and_result227[13]^and_result227[14]^and_result227[15]^and_result227[16]^and_result227[17]^and_result227[18]^and_result227[19]^and_result227[20]^and_result227[21]^and_result227[22]^and_result227[23]^and_result227[24]^and_result227[25]^and_result227[26]^and_result227[27]^and_result227[28]^and_result227[29]^and_result227[30]^and_result227[31]^and_result227[32]^and_result227[33]^and_result227[34]^and_result227[35]^and_result227[36]^and_result227[37]^and_result227[38]^and_result227[39]^and_result227[40]^and_result227[41]^and_result227[42]^and_result227[43]^and_result227[44]^and_result227[45]^and_result227[46]^and_result227[47]^and_result227[48]^and_result227[49]^and_result227[50]^and_result227[51]^and_result227[52]^and_result227[53]^and_result227[54]^and_result227[55]^and_result227[56]^and_result227[57]^and_result227[58]^and_result227[59]^and_result227[60]^and_result227[61]^and_result227[62]^and_result227[63]^and_result227[64]^and_result227[65]^and_result227[66]^and_result227[67]^and_result227[68]^and_result227[69]^and_result227[70]^and_result227[71]^and_result227[72]^and_result227[73]^and_result227[74]^and_result227[75]^and_result227[76]^and_result227[77]^and_result227[78]^and_result227[79]^and_result227[80]^and_result227[81]^and_result227[82]^and_result227[83]^and_result227[84]^and_result227[85]^and_result227[86]^and_result227[87]^and_result227[88]^and_result227[89]^and_result227[90]^and_result227[91]^and_result227[92]^and_result227[93]^and_result227[94]^and_result227[95]^and_result227[96]^and_result227[97]^and_result227[98]^and_result227[99]^and_result227[100]^and_result227[101]^and_result227[102]^and_result227[103]^and_result227[104]^and_result227[105]^and_result227[106]^and_result227[107]^and_result227[108]^and_result227[109]^and_result227[110]^and_result227[111]^and_result227[112]^and_result227[113]^and_result227[114]^and_result227[115]^and_result227[116]^and_result227[117]^and_result227[118]^and_result227[119]^and_result227[120]^and_result227[121]^and_result227[122]^and_result227[123]^and_result227[124]^and_result227[125]^and_result227[126]^and_result227[127]^and_result227[128]^and_result227[129]^and_result227[130]^and_result227[131]^and_result227[132]^and_result227[133]^and_result227[134]^and_result227[135]^and_result227[136]^and_result227[137]^and_result227[138]^and_result227[139]^and_result227[140]^and_result227[141]^and_result227[142]^and_result227[143]^and_result227[144]^and_result227[145]^and_result227[146]^and_result227[147]^and_result227[148]^and_result227[149]^and_result227[150]^and_result227[151]^and_result227[152]^and_result227[153]^and_result227[154]^and_result227[155]^and_result227[156]^and_result227[157]^and_result227[158]^and_result227[159]^and_result227[160]^and_result227[161]^and_result227[162]^and_result227[163]^and_result227[164]^and_result227[165]^and_result227[166]^and_result227[167]^and_result227[168]^and_result227[169]^and_result227[170]^and_result227[171]^and_result227[172]^and_result227[173]^and_result227[174]^and_result227[175]^and_result227[176]^and_result227[177]^and_result227[178]^and_result227[179]^and_result227[180]^and_result227[181]^and_result227[182]^and_result227[183]^and_result227[184]^and_result227[185]^and_result227[186]^and_result227[187]^and_result227[188]^and_result227[189]^and_result227[190]^and_result227[191]^and_result227[192]^and_result227[193]^and_result227[194]^and_result227[195]^and_result227[196]^and_result227[197]^and_result227[198]^and_result227[199]^and_result227[200]^and_result227[201]^and_result227[202]^and_result227[203]^and_result227[204]^and_result227[205]^and_result227[206]^and_result227[207]^and_result227[208]^and_result227[209]^and_result227[210]^and_result227[211]^and_result227[212]^and_result227[213]^and_result227[214]^and_result227[215]^and_result227[216]^and_result227[217]^and_result227[218]^and_result227[219]^and_result227[220]^and_result227[221]^and_result227[222]^and_result227[223]^and_result227[224]^and_result227[225]^and_result227[226]^and_result227[227]^and_result227[228]^and_result227[229]^and_result227[230]^and_result227[231]^and_result227[232]^and_result227[233]^and_result227[234]^and_result227[235]^and_result227[236]^and_result227[237]^and_result227[238]^and_result227[239]^and_result227[240]^and_result227[241]^and_result227[242]^and_result227[243]^and_result227[244]^and_result227[245]^and_result227[246]^and_result227[247]^and_result227[248]^and_result227[249]^and_result227[250]^and_result227[251]^and_result227[252]^and_result227[253]^and_result227[254];
assign key[228]=and_result228[0]^and_result228[1]^and_result228[2]^and_result228[3]^and_result228[4]^and_result228[5]^and_result228[6]^and_result228[7]^and_result228[8]^and_result228[9]^and_result228[10]^and_result228[11]^and_result228[12]^and_result228[13]^and_result228[14]^and_result228[15]^and_result228[16]^and_result228[17]^and_result228[18]^and_result228[19]^and_result228[20]^and_result228[21]^and_result228[22]^and_result228[23]^and_result228[24]^and_result228[25]^and_result228[26]^and_result228[27]^and_result228[28]^and_result228[29]^and_result228[30]^and_result228[31]^and_result228[32]^and_result228[33]^and_result228[34]^and_result228[35]^and_result228[36]^and_result228[37]^and_result228[38]^and_result228[39]^and_result228[40]^and_result228[41]^and_result228[42]^and_result228[43]^and_result228[44]^and_result228[45]^and_result228[46]^and_result228[47]^and_result228[48]^and_result228[49]^and_result228[50]^and_result228[51]^and_result228[52]^and_result228[53]^and_result228[54]^and_result228[55]^and_result228[56]^and_result228[57]^and_result228[58]^and_result228[59]^and_result228[60]^and_result228[61]^and_result228[62]^and_result228[63]^and_result228[64]^and_result228[65]^and_result228[66]^and_result228[67]^and_result228[68]^and_result228[69]^and_result228[70]^and_result228[71]^and_result228[72]^and_result228[73]^and_result228[74]^and_result228[75]^and_result228[76]^and_result228[77]^and_result228[78]^and_result228[79]^and_result228[80]^and_result228[81]^and_result228[82]^and_result228[83]^and_result228[84]^and_result228[85]^and_result228[86]^and_result228[87]^and_result228[88]^and_result228[89]^and_result228[90]^and_result228[91]^and_result228[92]^and_result228[93]^and_result228[94]^and_result228[95]^and_result228[96]^and_result228[97]^and_result228[98]^and_result228[99]^and_result228[100]^and_result228[101]^and_result228[102]^and_result228[103]^and_result228[104]^and_result228[105]^and_result228[106]^and_result228[107]^and_result228[108]^and_result228[109]^and_result228[110]^and_result228[111]^and_result228[112]^and_result228[113]^and_result228[114]^and_result228[115]^and_result228[116]^and_result228[117]^and_result228[118]^and_result228[119]^and_result228[120]^and_result228[121]^and_result228[122]^and_result228[123]^and_result228[124]^and_result228[125]^and_result228[126]^and_result228[127]^and_result228[128]^and_result228[129]^and_result228[130]^and_result228[131]^and_result228[132]^and_result228[133]^and_result228[134]^and_result228[135]^and_result228[136]^and_result228[137]^and_result228[138]^and_result228[139]^and_result228[140]^and_result228[141]^and_result228[142]^and_result228[143]^and_result228[144]^and_result228[145]^and_result228[146]^and_result228[147]^and_result228[148]^and_result228[149]^and_result228[150]^and_result228[151]^and_result228[152]^and_result228[153]^and_result228[154]^and_result228[155]^and_result228[156]^and_result228[157]^and_result228[158]^and_result228[159]^and_result228[160]^and_result228[161]^and_result228[162]^and_result228[163]^and_result228[164]^and_result228[165]^and_result228[166]^and_result228[167]^and_result228[168]^and_result228[169]^and_result228[170]^and_result228[171]^and_result228[172]^and_result228[173]^and_result228[174]^and_result228[175]^and_result228[176]^and_result228[177]^and_result228[178]^and_result228[179]^and_result228[180]^and_result228[181]^and_result228[182]^and_result228[183]^and_result228[184]^and_result228[185]^and_result228[186]^and_result228[187]^and_result228[188]^and_result228[189]^and_result228[190]^and_result228[191]^and_result228[192]^and_result228[193]^and_result228[194]^and_result228[195]^and_result228[196]^and_result228[197]^and_result228[198]^and_result228[199]^and_result228[200]^and_result228[201]^and_result228[202]^and_result228[203]^and_result228[204]^and_result228[205]^and_result228[206]^and_result228[207]^and_result228[208]^and_result228[209]^and_result228[210]^and_result228[211]^and_result228[212]^and_result228[213]^and_result228[214]^and_result228[215]^and_result228[216]^and_result228[217]^and_result228[218]^and_result228[219]^and_result228[220]^and_result228[221]^and_result228[222]^and_result228[223]^and_result228[224]^and_result228[225]^and_result228[226]^and_result228[227]^and_result228[228]^and_result228[229]^and_result228[230]^and_result228[231]^and_result228[232]^and_result228[233]^and_result228[234]^and_result228[235]^and_result228[236]^and_result228[237]^and_result228[238]^and_result228[239]^and_result228[240]^and_result228[241]^and_result228[242]^and_result228[243]^and_result228[244]^and_result228[245]^and_result228[246]^and_result228[247]^and_result228[248]^and_result228[249]^and_result228[250]^and_result228[251]^and_result228[252]^and_result228[253]^and_result228[254];
assign key[229]=and_result229[0]^and_result229[1]^and_result229[2]^and_result229[3]^and_result229[4]^and_result229[5]^and_result229[6]^and_result229[7]^and_result229[8]^and_result229[9]^and_result229[10]^and_result229[11]^and_result229[12]^and_result229[13]^and_result229[14]^and_result229[15]^and_result229[16]^and_result229[17]^and_result229[18]^and_result229[19]^and_result229[20]^and_result229[21]^and_result229[22]^and_result229[23]^and_result229[24]^and_result229[25]^and_result229[26]^and_result229[27]^and_result229[28]^and_result229[29]^and_result229[30]^and_result229[31]^and_result229[32]^and_result229[33]^and_result229[34]^and_result229[35]^and_result229[36]^and_result229[37]^and_result229[38]^and_result229[39]^and_result229[40]^and_result229[41]^and_result229[42]^and_result229[43]^and_result229[44]^and_result229[45]^and_result229[46]^and_result229[47]^and_result229[48]^and_result229[49]^and_result229[50]^and_result229[51]^and_result229[52]^and_result229[53]^and_result229[54]^and_result229[55]^and_result229[56]^and_result229[57]^and_result229[58]^and_result229[59]^and_result229[60]^and_result229[61]^and_result229[62]^and_result229[63]^and_result229[64]^and_result229[65]^and_result229[66]^and_result229[67]^and_result229[68]^and_result229[69]^and_result229[70]^and_result229[71]^and_result229[72]^and_result229[73]^and_result229[74]^and_result229[75]^and_result229[76]^and_result229[77]^and_result229[78]^and_result229[79]^and_result229[80]^and_result229[81]^and_result229[82]^and_result229[83]^and_result229[84]^and_result229[85]^and_result229[86]^and_result229[87]^and_result229[88]^and_result229[89]^and_result229[90]^and_result229[91]^and_result229[92]^and_result229[93]^and_result229[94]^and_result229[95]^and_result229[96]^and_result229[97]^and_result229[98]^and_result229[99]^and_result229[100]^and_result229[101]^and_result229[102]^and_result229[103]^and_result229[104]^and_result229[105]^and_result229[106]^and_result229[107]^and_result229[108]^and_result229[109]^and_result229[110]^and_result229[111]^and_result229[112]^and_result229[113]^and_result229[114]^and_result229[115]^and_result229[116]^and_result229[117]^and_result229[118]^and_result229[119]^and_result229[120]^and_result229[121]^and_result229[122]^and_result229[123]^and_result229[124]^and_result229[125]^and_result229[126]^and_result229[127]^and_result229[128]^and_result229[129]^and_result229[130]^and_result229[131]^and_result229[132]^and_result229[133]^and_result229[134]^and_result229[135]^and_result229[136]^and_result229[137]^and_result229[138]^and_result229[139]^and_result229[140]^and_result229[141]^and_result229[142]^and_result229[143]^and_result229[144]^and_result229[145]^and_result229[146]^and_result229[147]^and_result229[148]^and_result229[149]^and_result229[150]^and_result229[151]^and_result229[152]^and_result229[153]^and_result229[154]^and_result229[155]^and_result229[156]^and_result229[157]^and_result229[158]^and_result229[159]^and_result229[160]^and_result229[161]^and_result229[162]^and_result229[163]^and_result229[164]^and_result229[165]^and_result229[166]^and_result229[167]^and_result229[168]^and_result229[169]^and_result229[170]^and_result229[171]^and_result229[172]^and_result229[173]^and_result229[174]^and_result229[175]^and_result229[176]^and_result229[177]^and_result229[178]^and_result229[179]^and_result229[180]^and_result229[181]^and_result229[182]^and_result229[183]^and_result229[184]^and_result229[185]^and_result229[186]^and_result229[187]^and_result229[188]^and_result229[189]^and_result229[190]^and_result229[191]^and_result229[192]^and_result229[193]^and_result229[194]^and_result229[195]^and_result229[196]^and_result229[197]^and_result229[198]^and_result229[199]^and_result229[200]^and_result229[201]^and_result229[202]^and_result229[203]^and_result229[204]^and_result229[205]^and_result229[206]^and_result229[207]^and_result229[208]^and_result229[209]^and_result229[210]^and_result229[211]^and_result229[212]^and_result229[213]^and_result229[214]^and_result229[215]^and_result229[216]^and_result229[217]^and_result229[218]^and_result229[219]^and_result229[220]^and_result229[221]^and_result229[222]^and_result229[223]^and_result229[224]^and_result229[225]^and_result229[226]^and_result229[227]^and_result229[228]^and_result229[229]^and_result229[230]^and_result229[231]^and_result229[232]^and_result229[233]^and_result229[234]^and_result229[235]^and_result229[236]^and_result229[237]^and_result229[238]^and_result229[239]^and_result229[240]^and_result229[241]^and_result229[242]^and_result229[243]^and_result229[244]^and_result229[245]^and_result229[246]^and_result229[247]^and_result229[248]^and_result229[249]^and_result229[250]^and_result229[251]^and_result229[252]^and_result229[253]^and_result229[254];
assign key[230]=and_result230[0]^and_result230[1]^and_result230[2]^and_result230[3]^and_result230[4]^and_result230[5]^and_result230[6]^and_result230[7]^and_result230[8]^and_result230[9]^and_result230[10]^and_result230[11]^and_result230[12]^and_result230[13]^and_result230[14]^and_result230[15]^and_result230[16]^and_result230[17]^and_result230[18]^and_result230[19]^and_result230[20]^and_result230[21]^and_result230[22]^and_result230[23]^and_result230[24]^and_result230[25]^and_result230[26]^and_result230[27]^and_result230[28]^and_result230[29]^and_result230[30]^and_result230[31]^and_result230[32]^and_result230[33]^and_result230[34]^and_result230[35]^and_result230[36]^and_result230[37]^and_result230[38]^and_result230[39]^and_result230[40]^and_result230[41]^and_result230[42]^and_result230[43]^and_result230[44]^and_result230[45]^and_result230[46]^and_result230[47]^and_result230[48]^and_result230[49]^and_result230[50]^and_result230[51]^and_result230[52]^and_result230[53]^and_result230[54]^and_result230[55]^and_result230[56]^and_result230[57]^and_result230[58]^and_result230[59]^and_result230[60]^and_result230[61]^and_result230[62]^and_result230[63]^and_result230[64]^and_result230[65]^and_result230[66]^and_result230[67]^and_result230[68]^and_result230[69]^and_result230[70]^and_result230[71]^and_result230[72]^and_result230[73]^and_result230[74]^and_result230[75]^and_result230[76]^and_result230[77]^and_result230[78]^and_result230[79]^and_result230[80]^and_result230[81]^and_result230[82]^and_result230[83]^and_result230[84]^and_result230[85]^and_result230[86]^and_result230[87]^and_result230[88]^and_result230[89]^and_result230[90]^and_result230[91]^and_result230[92]^and_result230[93]^and_result230[94]^and_result230[95]^and_result230[96]^and_result230[97]^and_result230[98]^and_result230[99]^and_result230[100]^and_result230[101]^and_result230[102]^and_result230[103]^and_result230[104]^and_result230[105]^and_result230[106]^and_result230[107]^and_result230[108]^and_result230[109]^and_result230[110]^and_result230[111]^and_result230[112]^and_result230[113]^and_result230[114]^and_result230[115]^and_result230[116]^and_result230[117]^and_result230[118]^and_result230[119]^and_result230[120]^and_result230[121]^and_result230[122]^and_result230[123]^and_result230[124]^and_result230[125]^and_result230[126]^and_result230[127]^and_result230[128]^and_result230[129]^and_result230[130]^and_result230[131]^and_result230[132]^and_result230[133]^and_result230[134]^and_result230[135]^and_result230[136]^and_result230[137]^and_result230[138]^and_result230[139]^and_result230[140]^and_result230[141]^and_result230[142]^and_result230[143]^and_result230[144]^and_result230[145]^and_result230[146]^and_result230[147]^and_result230[148]^and_result230[149]^and_result230[150]^and_result230[151]^and_result230[152]^and_result230[153]^and_result230[154]^and_result230[155]^and_result230[156]^and_result230[157]^and_result230[158]^and_result230[159]^and_result230[160]^and_result230[161]^and_result230[162]^and_result230[163]^and_result230[164]^and_result230[165]^and_result230[166]^and_result230[167]^and_result230[168]^and_result230[169]^and_result230[170]^and_result230[171]^and_result230[172]^and_result230[173]^and_result230[174]^and_result230[175]^and_result230[176]^and_result230[177]^and_result230[178]^and_result230[179]^and_result230[180]^and_result230[181]^and_result230[182]^and_result230[183]^and_result230[184]^and_result230[185]^and_result230[186]^and_result230[187]^and_result230[188]^and_result230[189]^and_result230[190]^and_result230[191]^and_result230[192]^and_result230[193]^and_result230[194]^and_result230[195]^and_result230[196]^and_result230[197]^and_result230[198]^and_result230[199]^and_result230[200]^and_result230[201]^and_result230[202]^and_result230[203]^and_result230[204]^and_result230[205]^and_result230[206]^and_result230[207]^and_result230[208]^and_result230[209]^and_result230[210]^and_result230[211]^and_result230[212]^and_result230[213]^and_result230[214]^and_result230[215]^and_result230[216]^and_result230[217]^and_result230[218]^and_result230[219]^and_result230[220]^and_result230[221]^and_result230[222]^and_result230[223]^and_result230[224]^and_result230[225]^and_result230[226]^and_result230[227]^and_result230[228]^and_result230[229]^and_result230[230]^and_result230[231]^and_result230[232]^and_result230[233]^and_result230[234]^and_result230[235]^and_result230[236]^and_result230[237]^and_result230[238]^and_result230[239]^and_result230[240]^and_result230[241]^and_result230[242]^and_result230[243]^and_result230[244]^and_result230[245]^and_result230[246]^and_result230[247]^and_result230[248]^and_result230[249]^and_result230[250]^and_result230[251]^and_result230[252]^and_result230[253]^and_result230[254];
assign key[231]=and_result231[0]^and_result231[1]^and_result231[2]^and_result231[3]^and_result231[4]^and_result231[5]^and_result231[6]^and_result231[7]^and_result231[8]^and_result231[9]^and_result231[10]^and_result231[11]^and_result231[12]^and_result231[13]^and_result231[14]^and_result231[15]^and_result231[16]^and_result231[17]^and_result231[18]^and_result231[19]^and_result231[20]^and_result231[21]^and_result231[22]^and_result231[23]^and_result231[24]^and_result231[25]^and_result231[26]^and_result231[27]^and_result231[28]^and_result231[29]^and_result231[30]^and_result231[31]^and_result231[32]^and_result231[33]^and_result231[34]^and_result231[35]^and_result231[36]^and_result231[37]^and_result231[38]^and_result231[39]^and_result231[40]^and_result231[41]^and_result231[42]^and_result231[43]^and_result231[44]^and_result231[45]^and_result231[46]^and_result231[47]^and_result231[48]^and_result231[49]^and_result231[50]^and_result231[51]^and_result231[52]^and_result231[53]^and_result231[54]^and_result231[55]^and_result231[56]^and_result231[57]^and_result231[58]^and_result231[59]^and_result231[60]^and_result231[61]^and_result231[62]^and_result231[63]^and_result231[64]^and_result231[65]^and_result231[66]^and_result231[67]^and_result231[68]^and_result231[69]^and_result231[70]^and_result231[71]^and_result231[72]^and_result231[73]^and_result231[74]^and_result231[75]^and_result231[76]^and_result231[77]^and_result231[78]^and_result231[79]^and_result231[80]^and_result231[81]^and_result231[82]^and_result231[83]^and_result231[84]^and_result231[85]^and_result231[86]^and_result231[87]^and_result231[88]^and_result231[89]^and_result231[90]^and_result231[91]^and_result231[92]^and_result231[93]^and_result231[94]^and_result231[95]^and_result231[96]^and_result231[97]^and_result231[98]^and_result231[99]^and_result231[100]^and_result231[101]^and_result231[102]^and_result231[103]^and_result231[104]^and_result231[105]^and_result231[106]^and_result231[107]^and_result231[108]^and_result231[109]^and_result231[110]^and_result231[111]^and_result231[112]^and_result231[113]^and_result231[114]^and_result231[115]^and_result231[116]^and_result231[117]^and_result231[118]^and_result231[119]^and_result231[120]^and_result231[121]^and_result231[122]^and_result231[123]^and_result231[124]^and_result231[125]^and_result231[126]^and_result231[127]^and_result231[128]^and_result231[129]^and_result231[130]^and_result231[131]^and_result231[132]^and_result231[133]^and_result231[134]^and_result231[135]^and_result231[136]^and_result231[137]^and_result231[138]^and_result231[139]^and_result231[140]^and_result231[141]^and_result231[142]^and_result231[143]^and_result231[144]^and_result231[145]^and_result231[146]^and_result231[147]^and_result231[148]^and_result231[149]^and_result231[150]^and_result231[151]^and_result231[152]^and_result231[153]^and_result231[154]^and_result231[155]^and_result231[156]^and_result231[157]^and_result231[158]^and_result231[159]^and_result231[160]^and_result231[161]^and_result231[162]^and_result231[163]^and_result231[164]^and_result231[165]^and_result231[166]^and_result231[167]^and_result231[168]^and_result231[169]^and_result231[170]^and_result231[171]^and_result231[172]^and_result231[173]^and_result231[174]^and_result231[175]^and_result231[176]^and_result231[177]^and_result231[178]^and_result231[179]^and_result231[180]^and_result231[181]^and_result231[182]^and_result231[183]^and_result231[184]^and_result231[185]^and_result231[186]^and_result231[187]^and_result231[188]^and_result231[189]^and_result231[190]^and_result231[191]^and_result231[192]^and_result231[193]^and_result231[194]^and_result231[195]^and_result231[196]^and_result231[197]^and_result231[198]^and_result231[199]^and_result231[200]^and_result231[201]^and_result231[202]^and_result231[203]^and_result231[204]^and_result231[205]^and_result231[206]^and_result231[207]^and_result231[208]^and_result231[209]^and_result231[210]^and_result231[211]^and_result231[212]^and_result231[213]^and_result231[214]^and_result231[215]^and_result231[216]^and_result231[217]^and_result231[218]^and_result231[219]^and_result231[220]^and_result231[221]^and_result231[222]^and_result231[223]^and_result231[224]^and_result231[225]^and_result231[226]^and_result231[227]^and_result231[228]^and_result231[229]^and_result231[230]^and_result231[231]^and_result231[232]^and_result231[233]^and_result231[234]^and_result231[235]^and_result231[236]^and_result231[237]^and_result231[238]^and_result231[239]^and_result231[240]^and_result231[241]^and_result231[242]^and_result231[243]^and_result231[244]^and_result231[245]^and_result231[246]^and_result231[247]^and_result231[248]^and_result231[249]^and_result231[250]^and_result231[251]^and_result231[252]^and_result231[253]^and_result231[254];
assign key[232]=and_result232[0]^and_result232[1]^and_result232[2]^and_result232[3]^and_result232[4]^and_result232[5]^and_result232[6]^and_result232[7]^and_result232[8]^and_result232[9]^and_result232[10]^and_result232[11]^and_result232[12]^and_result232[13]^and_result232[14]^and_result232[15]^and_result232[16]^and_result232[17]^and_result232[18]^and_result232[19]^and_result232[20]^and_result232[21]^and_result232[22]^and_result232[23]^and_result232[24]^and_result232[25]^and_result232[26]^and_result232[27]^and_result232[28]^and_result232[29]^and_result232[30]^and_result232[31]^and_result232[32]^and_result232[33]^and_result232[34]^and_result232[35]^and_result232[36]^and_result232[37]^and_result232[38]^and_result232[39]^and_result232[40]^and_result232[41]^and_result232[42]^and_result232[43]^and_result232[44]^and_result232[45]^and_result232[46]^and_result232[47]^and_result232[48]^and_result232[49]^and_result232[50]^and_result232[51]^and_result232[52]^and_result232[53]^and_result232[54]^and_result232[55]^and_result232[56]^and_result232[57]^and_result232[58]^and_result232[59]^and_result232[60]^and_result232[61]^and_result232[62]^and_result232[63]^and_result232[64]^and_result232[65]^and_result232[66]^and_result232[67]^and_result232[68]^and_result232[69]^and_result232[70]^and_result232[71]^and_result232[72]^and_result232[73]^and_result232[74]^and_result232[75]^and_result232[76]^and_result232[77]^and_result232[78]^and_result232[79]^and_result232[80]^and_result232[81]^and_result232[82]^and_result232[83]^and_result232[84]^and_result232[85]^and_result232[86]^and_result232[87]^and_result232[88]^and_result232[89]^and_result232[90]^and_result232[91]^and_result232[92]^and_result232[93]^and_result232[94]^and_result232[95]^and_result232[96]^and_result232[97]^and_result232[98]^and_result232[99]^and_result232[100]^and_result232[101]^and_result232[102]^and_result232[103]^and_result232[104]^and_result232[105]^and_result232[106]^and_result232[107]^and_result232[108]^and_result232[109]^and_result232[110]^and_result232[111]^and_result232[112]^and_result232[113]^and_result232[114]^and_result232[115]^and_result232[116]^and_result232[117]^and_result232[118]^and_result232[119]^and_result232[120]^and_result232[121]^and_result232[122]^and_result232[123]^and_result232[124]^and_result232[125]^and_result232[126]^and_result232[127]^and_result232[128]^and_result232[129]^and_result232[130]^and_result232[131]^and_result232[132]^and_result232[133]^and_result232[134]^and_result232[135]^and_result232[136]^and_result232[137]^and_result232[138]^and_result232[139]^and_result232[140]^and_result232[141]^and_result232[142]^and_result232[143]^and_result232[144]^and_result232[145]^and_result232[146]^and_result232[147]^and_result232[148]^and_result232[149]^and_result232[150]^and_result232[151]^and_result232[152]^and_result232[153]^and_result232[154]^and_result232[155]^and_result232[156]^and_result232[157]^and_result232[158]^and_result232[159]^and_result232[160]^and_result232[161]^and_result232[162]^and_result232[163]^and_result232[164]^and_result232[165]^and_result232[166]^and_result232[167]^and_result232[168]^and_result232[169]^and_result232[170]^and_result232[171]^and_result232[172]^and_result232[173]^and_result232[174]^and_result232[175]^and_result232[176]^and_result232[177]^and_result232[178]^and_result232[179]^and_result232[180]^and_result232[181]^and_result232[182]^and_result232[183]^and_result232[184]^and_result232[185]^and_result232[186]^and_result232[187]^and_result232[188]^and_result232[189]^and_result232[190]^and_result232[191]^and_result232[192]^and_result232[193]^and_result232[194]^and_result232[195]^and_result232[196]^and_result232[197]^and_result232[198]^and_result232[199]^and_result232[200]^and_result232[201]^and_result232[202]^and_result232[203]^and_result232[204]^and_result232[205]^and_result232[206]^and_result232[207]^and_result232[208]^and_result232[209]^and_result232[210]^and_result232[211]^and_result232[212]^and_result232[213]^and_result232[214]^and_result232[215]^and_result232[216]^and_result232[217]^and_result232[218]^and_result232[219]^and_result232[220]^and_result232[221]^and_result232[222]^and_result232[223]^and_result232[224]^and_result232[225]^and_result232[226]^and_result232[227]^and_result232[228]^and_result232[229]^and_result232[230]^and_result232[231]^and_result232[232]^and_result232[233]^and_result232[234]^and_result232[235]^and_result232[236]^and_result232[237]^and_result232[238]^and_result232[239]^and_result232[240]^and_result232[241]^and_result232[242]^and_result232[243]^and_result232[244]^and_result232[245]^and_result232[246]^and_result232[247]^and_result232[248]^and_result232[249]^and_result232[250]^and_result232[251]^and_result232[252]^and_result232[253]^and_result232[254];
assign key[233]=and_result233[0]^and_result233[1]^and_result233[2]^and_result233[3]^and_result233[4]^and_result233[5]^and_result233[6]^and_result233[7]^and_result233[8]^and_result233[9]^and_result233[10]^and_result233[11]^and_result233[12]^and_result233[13]^and_result233[14]^and_result233[15]^and_result233[16]^and_result233[17]^and_result233[18]^and_result233[19]^and_result233[20]^and_result233[21]^and_result233[22]^and_result233[23]^and_result233[24]^and_result233[25]^and_result233[26]^and_result233[27]^and_result233[28]^and_result233[29]^and_result233[30]^and_result233[31]^and_result233[32]^and_result233[33]^and_result233[34]^and_result233[35]^and_result233[36]^and_result233[37]^and_result233[38]^and_result233[39]^and_result233[40]^and_result233[41]^and_result233[42]^and_result233[43]^and_result233[44]^and_result233[45]^and_result233[46]^and_result233[47]^and_result233[48]^and_result233[49]^and_result233[50]^and_result233[51]^and_result233[52]^and_result233[53]^and_result233[54]^and_result233[55]^and_result233[56]^and_result233[57]^and_result233[58]^and_result233[59]^and_result233[60]^and_result233[61]^and_result233[62]^and_result233[63]^and_result233[64]^and_result233[65]^and_result233[66]^and_result233[67]^and_result233[68]^and_result233[69]^and_result233[70]^and_result233[71]^and_result233[72]^and_result233[73]^and_result233[74]^and_result233[75]^and_result233[76]^and_result233[77]^and_result233[78]^and_result233[79]^and_result233[80]^and_result233[81]^and_result233[82]^and_result233[83]^and_result233[84]^and_result233[85]^and_result233[86]^and_result233[87]^and_result233[88]^and_result233[89]^and_result233[90]^and_result233[91]^and_result233[92]^and_result233[93]^and_result233[94]^and_result233[95]^and_result233[96]^and_result233[97]^and_result233[98]^and_result233[99]^and_result233[100]^and_result233[101]^and_result233[102]^and_result233[103]^and_result233[104]^and_result233[105]^and_result233[106]^and_result233[107]^and_result233[108]^and_result233[109]^and_result233[110]^and_result233[111]^and_result233[112]^and_result233[113]^and_result233[114]^and_result233[115]^and_result233[116]^and_result233[117]^and_result233[118]^and_result233[119]^and_result233[120]^and_result233[121]^and_result233[122]^and_result233[123]^and_result233[124]^and_result233[125]^and_result233[126]^and_result233[127]^and_result233[128]^and_result233[129]^and_result233[130]^and_result233[131]^and_result233[132]^and_result233[133]^and_result233[134]^and_result233[135]^and_result233[136]^and_result233[137]^and_result233[138]^and_result233[139]^and_result233[140]^and_result233[141]^and_result233[142]^and_result233[143]^and_result233[144]^and_result233[145]^and_result233[146]^and_result233[147]^and_result233[148]^and_result233[149]^and_result233[150]^and_result233[151]^and_result233[152]^and_result233[153]^and_result233[154]^and_result233[155]^and_result233[156]^and_result233[157]^and_result233[158]^and_result233[159]^and_result233[160]^and_result233[161]^and_result233[162]^and_result233[163]^and_result233[164]^and_result233[165]^and_result233[166]^and_result233[167]^and_result233[168]^and_result233[169]^and_result233[170]^and_result233[171]^and_result233[172]^and_result233[173]^and_result233[174]^and_result233[175]^and_result233[176]^and_result233[177]^and_result233[178]^and_result233[179]^and_result233[180]^and_result233[181]^and_result233[182]^and_result233[183]^and_result233[184]^and_result233[185]^and_result233[186]^and_result233[187]^and_result233[188]^and_result233[189]^and_result233[190]^and_result233[191]^and_result233[192]^and_result233[193]^and_result233[194]^and_result233[195]^and_result233[196]^and_result233[197]^and_result233[198]^and_result233[199]^and_result233[200]^and_result233[201]^and_result233[202]^and_result233[203]^and_result233[204]^and_result233[205]^and_result233[206]^and_result233[207]^and_result233[208]^and_result233[209]^and_result233[210]^and_result233[211]^and_result233[212]^and_result233[213]^and_result233[214]^and_result233[215]^and_result233[216]^and_result233[217]^and_result233[218]^and_result233[219]^and_result233[220]^and_result233[221]^and_result233[222]^and_result233[223]^and_result233[224]^and_result233[225]^and_result233[226]^and_result233[227]^and_result233[228]^and_result233[229]^and_result233[230]^and_result233[231]^and_result233[232]^and_result233[233]^and_result233[234]^and_result233[235]^and_result233[236]^and_result233[237]^and_result233[238]^and_result233[239]^and_result233[240]^and_result233[241]^and_result233[242]^and_result233[243]^and_result233[244]^and_result233[245]^and_result233[246]^and_result233[247]^and_result233[248]^and_result233[249]^and_result233[250]^and_result233[251]^and_result233[252]^and_result233[253]^and_result233[254];
assign key[234]=and_result234[0]^and_result234[1]^and_result234[2]^and_result234[3]^and_result234[4]^and_result234[5]^and_result234[6]^and_result234[7]^and_result234[8]^and_result234[9]^and_result234[10]^and_result234[11]^and_result234[12]^and_result234[13]^and_result234[14]^and_result234[15]^and_result234[16]^and_result234[17]^and_result234[18]^and_result234[19]^and_result234[20]^and_result234[21]^and_result234[22]^and_result234[23]^and_result234[24]^and_result234[25]^and_result234[26]^and_result234[27]^and_result234[28]^and_result234[29]^and_result234[30]^and_result234[31]^and_result234[32]^and_result234[33]^and_result234[34]^and_result234[35]^and_result234[36]^and_result234[37]^and_result234[38]^and_result234[39]^and_result234[40]^and_result234[41]^and_result234[42]^and_result234[43]^and_result234[44]^and_result234[45]^and_result234[46]^and_result234[47]^and_result234[48]^and_result234[49]^and_result234[50]^and_result234[51]^and_result234[52]^and_result234[53]^and_result234[54]^and_result234[55]^and_result234[56]^and_result234[57]^and_result234[58]^and_result234[59]^and_result234[60]^and_result234[61]^and_result234[62]^and_result234[63]^and_result234[64]^and_result234[65]^and_result234[66]^and_result234[67]^and_result234[68]^and_result234[69]^and_result234[70]^and_result234[71]^and_result234[72]^and_result234[73]^and_result234[74]^and_result234[75]^and_result234[76]^and_result234[77]^and_result234[78]^and_result234[79]^and_result234[80]^and_result234[81]^and_result234[82]^and_result234[83]^and_result234[84]^and_result234[85]^and_result234[86]^and_result234[87]^and_result234[88]^and_result234[89]^and_result234[90]^and_result234[91]^and_result234[92]^and_result234[93]^and_result234[94]^and_result234[95]^and_result234[96]^and_result234[97]^and_result234[98]^and_result234[99]^and_result234[100]^and_result234[101]^and_result234[102]^and_result234[103]^and_result234[104]^and_result234[105]^and_result234[106]^and_result234[107]^and_result234[108]^and_result234[109]^and_result234[110]^and_result234[111]^and_result234[112]^and_result234[113]^and_result234[114]^and_result234[115]^and_result234[116]^and_result234[117]^and_result234[118]^and_result234[119]^and_result234[120]^and_result234[121]^and_result234[122]^and_result234[123]^and_result234[124]^and_result234[125]^and_result234[126]^and_result234[127]^and_result234[128]^and_result234[129]^and_result234[130]^and_result234[131]^and_result234[132]^and_result234[133]^and_result234[134]^and_result234[135]^and_result234[136]^and_result234[137]^and_result234[138]^and_result234[139]^and_result234[140]^and_result234[141]^and_result234[142]^and_result234[143]^and_result234[144]^and_result234[145]^and_result234[146]^and_result234[147]^and_result234[148]^and_result234[149]^and_result234[150]^and_result234[151]^and_result234[152]^and_result234[153]^and_result234[154]^and_result234[155]^and_result234[156]^and_result234[157]^and_result234[158]^and_result234[159]^and_result234[160]^and_result234[161]^and_result234[162]^and_result234[163]^and_result234[164]^and_result234[165]^and_result234[166]^and_result234[167]^and_result234[168]^and_result234[169]^and_result234[170]^and_result234[171]^and_result234[172]^and_result234[173]^and_result234[174]^and_result234[175]^and_result234[176]^and_result234[177]^and_result234[178]^and_result234[179]^and_result234[180]^and_result234[181]^and_result234[182]^and_result234[183]^and_result234[184]^and_result234[185]^and_result234[186]^and_result234[187]^and_result234[188]^and_result234[189]^and_result234[190]^and_result234[191]^and_result234[192]^and_result234[193]^and_result234[194]^and_result234[195]^and_result234[196]^and_result234[197]^and_result234[198]^and_result234[199]^and_result234[200]^and_result234[201]^and_result234[202]^and_result234[203]^and_result234[204]^and_result234[205]^and_result234[206]^and_result234[207]^and_result234[208]^and_result234[209]^and_result234[210]^and_result234[211]^and_result234[212]^and_result234[213]^and_result234[214]^and_result234[215]^and_result234[216]^and_result234[217]^and_result234[218]^and_result234[219]^and_result234[220]^and_result234[221]^and_result234[222]^and_result234[223]^and_result234[224]^and_result234[225]^and_result234[226]^and_result234[227]^and_result234[228]^and_result234[229]^and_result234[230]^and_result234[231]^and_result234[232]^and_result234[233]^and_result234[234]^and_result234[235]^and_result234[236]^and_result234[237]^and_result234[238]^and_result234[239]^and_result234[240]^and_result234[241]^and_result234[242]^and_result234[243]^and_result234[244]^and_result234[245]^and_result234[246]^and_result234[247]^and_result234[248]^and_result234[249]^and_result234[250]^and_result234[251]^and_result234[252]^and_result234[253]^and_result234[254];
assign key[235]=and_result235[0]^and_result235[1]^and_result235[2]^and_result235[3]^and_result235[4]^and_result235[5]^and_result235[6]^and_result235[7]^and_result235[8]^and_result235[9]^and_result235[10]^and_result235[11]^and_result235[12]^and_result235[13]^and_result235[14]^and_result235[15]^and_result235[16]^and_result235[17]^and_result235[18]^and_result235[19]^and_result235[20]^and_result235[21]^and_result235[22]^and_result235[23]^and_result235[24]^and_result235[25]^and_result235[26]^and_result235[27]^and_result235[28]^and_result235[29]^and_result235[30]^and_result235[31]^and_result235[32]^and_result235[33]^and_result235[34]^and_result235[35]^and_result235[36]^and_result235[37]^and_result235[38]^and_result235[39]^and_result235[40]^and_result235[41]^and_result235[42]^and_result235[43]^and_result235[44]^and_result235[45]^and_result235[46]^and_result235[47]^and_result235[48]^and_result235[49]^and_result235[50]^and_result235[51]^and_result235[52]^and_result235[53]^and_result235[54]^and_result235[55]^and_result235[56]^and_result235[57]^and_result235[58]^and_result235[59]^and_result235[60]^and_result235[61]^and_result235[62]^and_result235[63]^and_result235[64]^and_result235[65]^and_result235[66]^and_result235[67]^and_result235[68]^and_result235[69]^and_result235[70]^and_result235[71]^and_result235[72]^and_result235[73]^and_result235[74]^and_result235[75]^and_result235[76]^and_result235[77]^and_result235[78]^and_result235[79]^and_result235[80]^and_result235[81]^and_result235[82]^and_result235[83]^and_result235[84]^and_result235[85]^and_result235[86]^and_result235[87]^and_result235[88]^and_result235[89]^and_result235[90]^and_result235[91]^and_result235[92]^and_result235[93]^and_result235[94]^and_result235[95]^and_result235[96]^and_result235[97]^and_result235[98]^and_result235[99]^and_result235[100]^and_result235[101]^and_result235[102]^and_result235[103]^and_result235[104]^and_result235[105]^and_result235[106]^and_result235[107]^and_result235[108]^and_result235[109]^and_result235[110]^and_result235[111]^and_result235[112]^and_result235[113]^and_result235[114]^and_result235[115]^and_result235[116]^and_result235[117]^and_result235[118]^and_result235[119]^and_result235[120]^and_result235[121]^and_result235[122]^and_result235[123]^and_result235[124]^and_result235[125]^and_result235[126]^and_result235[127]^and_result235[128]^and_result235[129]^and_result235[130]^and_result235[131]^and_result235[132]^and_result235[133]^and_result235[134]^and_result235[135]^and_result235[136]^and_result235[137]^and_result235[138]^and_result235[139]^and_result235[140]^and_result235[141]^and_result235[142]^and_result235[143]^and_result235[144]^and_result235[145]^and_result235[146]^and_result235[147]^and_result235[148]^and_result235[149]^and_result235[150]^and_result235[151]^and_result235[152]^and_result235[153]^and_result235[154]^and_result235[155]^and_result235[156]^and_result235[157]^and_result235[158]^and_result235[159]^and_result235[160]^and_result235[161]^and_result235[162]^and_result235[163]^and_result235[164]^and_result235[165]^and_result235[166]^and_result235[167]^and_result235[168]^and_result235[169]^and_result235[170]^and_result235[171]^and_result235[172]^and_result235[173]^and_result235[174]^and_result235[175]^and_result235[176]^and_result235[177]^and_result235[178]^and_result235[179]^and_result235[180]^and_result235[181]^and_result235[182]^and_result235[183]^and_result235[184]^and_result235[185]^and_result235[186]^and_result235[187]^and_result235[188]^and_result235[189]^and_result235[190]^and_result235[191]^and_result235[192]^and_result235[193]^and_result235[194]^and_result235[195]^and_result235[196]^and_result235[197]^and_result235[198]^and_result235[199]^and_result235[200]^and_result235[201]^and_result235[202]^and_result235[203]^and_result235[204]^and_result235[205]^and_result235[206]^and_result235[207]^and_result235[208]^and_result235[209]^and_result235[210]^and_result235[211]^and_result235[212]^and_result235[213]^and_result235[214]^and_result235[215]^and_result235[216]^and_result235[217]^and_result235[218]^and_result235[219]^and_result235[220]^and_result235[221]^and_result235[222]^and_result235[223]^and_result235[224]^and_result235[225]^and_result235[226]^and_result235[227]^and_result235[228]^and_result235[229]^and_result235[230]^and_result235[231]^and_result235[232]^and_result235[233]^and_result235[234]^and_result235[235]^and_result235[236]^and_result235[237]^and_result235[238]^and_result235[239]^and_result235[240]^and_result235[241]^and_result235[242]^and_result235[243]^and_result235[244]^and_result235[245]^and_result235[246]^and_result235[247]^and_result235[248]^and_result235[249]^and_result235[250]^and_result235[251]^and_result235[252]^and_result235[253]^and_result235[254];
assign key[236]=and_result236[0]^and_result236[1]^and_result236[2]^and_result236[3]^and_result236[4]^and_result236[5]^and_result236[6]^and_result236[7]^and_result236[8]^and_result236[9]^and_result236[10]^and_result236[11]^and_result236[12]^and_result236[13]^and_result236[14]^and_result236[15]^and_result236[16]^and_result236[17]^and_result236[18]^and_result236[19]^and_result236[20]^and_result236[21]^and_result236[22]^and_result236[23]^and_result236[24]^and_result236[25]^and_result236[26]^and_result236[27]^and_result236[28]^and_result236[29]^and_result236[30]^and_result236[31]^and_result236[32]^and_result236[33]^and_result236[34]^and_result236[35]^and_result236[36]^and_result236[37]^and_result236[38]^and_result236[39]^and_result236[40]^and_result236[41]^and_result236[42]^and_result236[43]^and_result236[44]^and_result236[45]^and_result236[46]^and_result236[47]^and_result236[48]^and_result236[49]^and_result236[50]^and_result236[51]^and_result236[52]^and_result236[53]^and_result236[54]^and_result236[55]^and_result236[56]^and_result236[57]^and_result236[58]^and_result236[59]^and_result236[60]^and_result236[61]^and_result236[62]^and_result236[63]^and_result236[64]^and_result236[65]^and_result236[66]^and_result236[67]^and_result236[68]^and_result236[69]^and_result236[70]^and_result236[71]^and_result236[72]^and_result236[73]^and_result236[74]^and_result236[75]^and_result236[76]^and_result236[77]^and_result236[78]^and_result236[79]^and_result236[80]^and_result236[81]^and_result236[82]^and_result236[83]^and_result236[84]^and_result236[85]^and_result236[86]^and_result236[87]^and_result236[88]^and_result236[89]^and_result236[90]^and_result236[91]^and_result236[92]^and_result236[93]^and_result236[94]^and_result236[95]^and_result236[96]^and_result236[97]^and_result236[98]^and_result236[99]^and_result236[100]^and_result236[101]^and_result236[102]^and_result236[103]^and_result236[104]^and_result236[105]^and_result236[106]^and_result236[107]^and_result236[108]^and_result236[109]^and_result236[110]^and_result236[111]^and_result236[112]^and_result236[113]^and_result236[114]^and_result236[115]^and_result236[116]^and_result236[117]^and_result236[118]^and_result236[119]^and_result236[120]^and_result236[121]^and_result236[122]^and_result236[123]^and_result236[124]^and_result236[125]^and_result236[126]^and_result236[127]^and_result236[128]^and_result236[129]^and_result236[130]^and_result236[131]^and_result236[132]^and_result236[133]^and_result236[134]^and_result236[135]^and_result236[136]^and_result236[137]^and_result236[138]^and_result236[139]^and_result236[140]^and_result236[141]^and_result236[142]^and_result236[143]^and_result236[144]^and_result236[145]^and_result236[146]^and_result236[147]^and_result236[148]^and_result236[149]^and_result236[150]^and_result236[151]^and_result236[152]^and_result236[153]^and_result236[154]^and_result236[155]^and_result236[156]^and_result236[157]^and_result236[158]^and_result236[159]^and_result236[160]^and_result236[161]^and_result236[162]^and_result236[163]^and_result236[164]^and_result236[165]^and_result236[166]^and_result236[167]^and_result236[168]^and_result236[169]^and_result236[170]^and_result236[171]^and_result236[172]^and_result236[173]^and_result236[174]^and_result236[175]^and_result236[176]^and_result236[177]^and_result236[178]^and_result236[179]^and_result236[180]^and_result236[181]^and_result236[182]^and_result236[183]^and_result236[184]^and_result236[185]^and_result236[186]^and_result236[187]^and_result236[188]^and_result236[189]^and_result236[190]^and_result236[191]^and_result236[192]^and_result236[193]^and_result236[194]^and_result236[195]^and_result236[196]^and_result236[197]^and_result236[198]^and_result236[199]^and_result236[200]^and_result236[201]^and_result236[202]^and_result236[203]^and_result236[204]^and_result236[205]^and_result236[206]^and_result236[207]^and_result236[208]^and_result236[209]^and_result236[210]^and_result236[211]^and_result236[212]^and_result236[213]^and_result236[214]^and_result236[215]^and_result236[216]^and_result236[217]^and_result236[218]^and_result236[219]^and_result236[220]^and_result236[221]^and_result236[222]^and_result236[223]^and_result236[224]^and_result236[225]^and_result236[226]^and_result236[227]^and_result236[228]^and_result236[229]^and_result236[230]^and_result236[231]^and_result236[232]^and_result236[233]^and_result236[234]^and_result236[235]^and_result236[236]^and_result236[237]^and_result236[238]^and_result236[239]^and_result236[240]^and_result236[241]^and_result236[242]^and_result236[243]^and_result236[244]^and_result236[245]^and_result236[246]^and_result236[247]^and_result236[248]^and_result236[249]^and_result236[250]^and_result236[251]^and_result236[252]^and_result236[253]^and_result236[254];
assign key[237]=and_result237[0]^and_result237[1]^and_result237[2]^and_result237[3]^and_result237[4]^and_result237[5]^and_result237[6]^and_result237[7]^and_result237[8]^and_result237[9]^and_result237[10]^and_result237[11]^and_result237[12]^and_result237[13]^and_result237[14]^and_result237[15]^and_result237[16]^and_result237[17]^and_result237[18]^and_result237[19]^and_result237[20]^and_result237[21]^and_result237[22]^and_result237[23]^and_result237[24]^and_result237[25]^and_result237[26]^and_result237[27]^and_result237[28]^and_result237[29]^and_result237[30]^and_result237[31]^and_result237[32]^and_result237[33]^and_result237[34]^and_result237[35]^and_result237[36]^and_result237[37]^and_result237[38]^and_result237[39]^and_result237[40]^and_result237[41]^and_result237[42]^and_result237[43]^and_result237[44]^and_result237[45]^and_result237[46]^and_result237[47]^and_result237[48]^and_result237[49]^and_result237[50]^and_result237[51]^and_result237[52]^and_result237[53]^and_result237[54]^and_result237[55]^and_result237[56]^and_result237[57]^and_result237[58]^and_result237[59]^and_result237[60]^and_result237[61]^and_result237[62]^and_result237[63]^and_result237[64]^and_result237[65]^and_result237[66]^and_result237[67]^and_result237[68]^and_result237[69]^and_result237[70]^and_result237[71]^and_result237[72]^and_result237[73]^and_result237[74]^and_result237[75]^and_result237[76]^and_result237[77]^and_result237[78]^and_result237[79]^and_result237[80]^and_result237[81]^and_result237[82]^and_result237[83]^and_result237[84]^and_result237[85]^and_result237[86]^and_result237[87]^and_result237[88]^and_result237[89]^and_result237[90]^and_result237[91]^and_result237[92]^and_result237[93]^and_result237[94]^and_result237[95]^and_result237[96]^and_result237[97]^and_result237[98]^and_result237[99]^and_result237[100]^and_result237[101]^and_result237[102]^and_result237[103]^and_result237[104]^and_result237[105]^and_result237[106]^and_result237[107]^and_result237[108]^and_result237[109]^and_result237[110]^and_result237[111]^and_result237[112]^and_result237[113]^and_result237[114]^and_result237[115]^and_result237[116]^and_result237[117]^and_result237[118]^and_result237[119]^and_result237[120]^and_result237[121]^and_result237[122]^and_result237[123]^and_result237[124]^and_result237[125]^and_result237[126]^and_result237[127]^and_result237[128]^and_result237[129]^and_result237[130]^and_result237[131]^and_result237[132]^and_result237[133]^and_result237[134]^and_result237[135]^and_result237[136]^and_result237[137]^and_result237[138]^and_result237[139]^and_result237[140]^and_result237[141]^and_result237[142]^and_result237[143]^and_result237[144]^and_result237[145]^and_result237[146]^and_result237[147]^and_result237[148]^and_result237[149]^and_result237[150]^and_result237[151]^and_result237[152]^and_result237[153]^and_result237[154]^and_result237[155]^and_result237[156]^and_result237[157]^and_result237[158]^and_result237[159]^and_result237[160]^and_result237[161]^and_result237[162]^and_result237[163]^and_result237[164]^and_result237[165]^and_result237[166]^and_result237[167]^and_result237[168]^and_result237[169]^and_result237[170]^and_result237[171]^and_result237[172]^and_result237[173]^and_result237[174]^and_result237[175]^and_result237[176]^and_result237[177]^and_result237[178]^and_result237[179]^and_result237[180]^and_result237[181]^and_result237[182]^and_result237[183]^and_result237[184]^and_result237[185]^and_result237[186]^and_result237[187]^and_result237[188]^and_result237[189]^and_result237[190]^and_result237[191]^and_result237[192]^and_result237[193]^and_result237[194]^and_result237[195]^and_result237[196]^and_result237[197]^and_result237[198]^and_result237[199]^and_result237[200]^and_result237[201]^and_result237[202]^and_result237[203]^and_result237[204]^and_result237[205]^and_result237[206]^and_result237[207]^and_result237[208]^and_result237[209]^and_result237[210]^and_result237[211]^and_result237[212]^and_result237[213]^and_result237[214]^and_result237[215]^and_result237[216]^and_result237[217]^and_result237[218]^and_result237[219]^and_result237[220]^and_result237[221]^and_result237[222]^and_result237[223]^and_result237[224]^and_result237[225]^and_result237[226]^and_result237[227]^and_result237[228]^and_result237[229]^and_result237[230]^and_result237[231]^and_result237[232]^and_result237[233]^and_result237[234]^and_result237[235]^and_result237[236]^and_result237[237]^and_result237[238]^and_result237[239]^and_result237[240]^and_result237[241]^and_result237[242]^and_result237[243]^and_result237[244]^and_result237[245]^and_result237[246]^and_result237[247]^and_result237[248]^and_result237[249]^and_result237[250]^and_result237[251]^and_result237[252]^and_result237[253]^and_result237[254];
assign key[238]=and_result238[0]^and_result238[1]^and_result238[2]^and_result238[3]^and_result238[4]^and_result238[5]^and_result238[6]^and_result238[7]^and_result238[8]^and_result238[9]^and_result238[10]^and_result238[11]^and_result238[12]^and_result238[13]^and_result238[14]^and_result238[15]^and_result238[16]^and_result238[17]^and_result238[18]^and_result238[19]^and_result238[20]^and_result238[21]^and_result238[22]^and_result238[23]^and_result238[24]^and_result238[25]^and_result238[26]^and_result238[27]^and_result238[28]^and_result238[29]^and_result238[30]^and_result238[31]^and_result238[32]^and_result238[33]^and_result238[34]^and_result238[35]^and_result238[36]^and_result238[37]^and_result238[38]^and_result238[39]^and_result238[40]^and_result238[41]^and_result238[42]^and_result238[43]^and_result238[44]^and_result238[45]^and_result238[46]^and_result238[47]^and_result238[48]^and_result238[49]^and_result238[50]^and_result238[51]^and_result238[52]^and_result238[53]^and_result238[54]^and_result238[55]^and_result238[56]^and_result238[57]^and_result238[58]^and_result238[59]^and_result238[60]^and_result238[61]^and_result238[62]^and_result238[63]^and_result238[64]^and_result238[65]^and_result238[66]^and_result238[67]^and_result238[68]^and_result238[69]^and_result238[70]^and_result238[71]^and_result238[72]^and_result238[73]^and_result238[74]^and_result238[75]^and_result238[76]^and_result238[77]^and_result238[78]^and_result238[79]^and_result238[80]^and_result238[81]^and_result238[82]^and_result238[83]^and_result238[84]^and_result238[85]^and_result238[86]^and_result238[87]^and_result238[88]^and_result238[89]^and_result238[90]^and_result238[91]^and_result238[92]^and_result238[93]^and_result238[94]^and_result238[95]^and_result238[96]^and_result238[97]^and_result238[98]^and_result238[99]^and_result238[100]^and_result238[101]^and_result238[102]^and_result238[103]^and_result238[104]^and_result238[105]^and_result238[106]^and_result238[107]^and_result238[108]^and_result238[109]^and_result238[110]^and_result238[111]^and_result238[112]^and_result238[113]^and_result238[114]^and_result238[115]^and_result238[116]^and_result238[117]^and_result238[118]^and_result238[119]^and_result238[120]^and_result238[121]^and_result238[122]^and_result238[123]^and_result238[124]^and_result238[125]^and_result238[126]^and_result238[127]^and_result238[128]^and_result238[129]^and_result238[130]^and_result238[131]^and_result238[132]^and_result238[133]^and_result238[134]^and_result238[135]^and_result238[136]^and_result238[137]^and_result238[138]^and_result238[139]^and_result238[140]^and_result238[141]^and_result238[142]^and_result238[143]^and_result238[144]^and_result238[145]^and_result238[146]^and_result238[147]^and_result238[148]^and_result238[149]^and_result238[150]^and_result238[151]^and_result238[152]^and_result238[153]^and_result238[154]^and_result238[155]^and_result238[156]^and_result238[157]^and_result238[158]^and_result238[159]^and_result238[160]^and_result238[161]^and_result238[162]^and_result238[163]^and_result238[164]^and_result238[165]^and_result238[166]^and_result238[167]^and_result238[168]^and_result238[169]^and_result238[170]^and_result238[171]^and_result238[172]^and_result238[173]^and_result238[174]^and_result238[175]^and_result238[176]^and_result238[177]^and_result238[178]^and_result238[179]^and_result238[180]^and_result238[181]^and_result238[182]^and_result238[183]^and_result238[184]^and_result238[185]^and_result238[186]^and_result238[187]^and_result238[188]^and_result238[189]^and_result238[190]^and_result238[191]^and_result238[192]^and_result238[193]^and_result238[194]^and_result238[195]^and_result238[196]^and_result238[197]^and_result238[198]^and_result238[199]^and_result238[200]^and_result238[201]^and_result238[202]^and_result238[203]^and_result238[204]^and_result238[205]^and_result238[206]^and_result238[207]^and_result238[208]^and_result238[209]^and_result238[210]^and_result238[211]^and_result238[212]^and_result238[213]^and_result238[214]^and_result238[215]^and_result238[216]^and_result238[217]^and_result238[218]^and_result238[219]^and_result238[220]^and_result238[221]^and_result238[222]^and_result238[223]^and_result238[224]^and_result238[225]^and_result238[226]^and_result238[227]^and_result238[228]^and_result238[229]^and_result238[230]^and_result238[231]^and_result238[232]^and_result238[233]^and_result238[234]^and_result238[235]^and_result238[236]^and_result238[237]^and_result238[238]^and_result238[239]^and_result238[240]^and_result238[241]^and_result238[242]^and_result238[243]^and_result238[244]^and_result238[245]^and_result238[246]^and_result238[247]^and_result238[248]^and_result238[249]^and_result238[250]^and_result238[251]^and_result238[252]^and_result238[253]^and_result238[254];
assign key[239]=and_result239[0]^and_result239[1]^and_result239[2]^and_result239[3]^and_result239[4]^and_result239[5]^and_result239[6]^and_result239[7]^and_result239[8]^and_result239[9]^and_result239[10]^and_result239[11]^and_result239[12]^and_result239[13]^and_result239[14]^and_result239[15]^and_result239[16]^and_result239[17]^and_result239[18]^and_result239[19]^and_result239[20]^and_result239[21]^and_result239[22]^and_result239[23]^and_result239[24]^and_result239[25]^and_result239[26]^and_result239[27]^and_result239[28]^and_result239[29]^and_result239[30]^and_result239[31]^and_result239[32]^and_result239[33]^and_result239[34]^and_result239[35]^and_result239[36]^and_result239[37]^and_result239[38]^and_result239[39]^and_result239[40]^and_result239[41]^and_result239[42]^and_result239[43]^and_result239[44]^and_result239[45]^and_result239[46]^and_result239[47]^and_result239[48]^and_result239[49]^and_result239[50]^and_result239[51]^and_result239[52]^and_result239[53]^and_result239[54]^and_result239[55]^and_result239[56]^and_result239[57]^and_result239[58]^and_result239[59]^and_result239[60]^and_result239[61]^and_result239[62]^and_result239[63]^and_result239[64]^and_result239[65]^and_result239[66]^and_result239[67]^and_result239[68]^and_result239[69]^and_result239[70]^and_result239[71]^and_result239[72]^and_result239[73]^and_result239[74]^and_result239[75]^and_result239[76]^and_result239[77]^and_result239[78]^and_result239[79]^and_result239[80]^and_result239[81]^and_result239[82]^and_result239[83]^and_result239[84]^and_result239[85]^and_result239[86]^and_result239[87]^and_result239[88]^and_result239[89]^and_result239[90]^and_result239[91]^and_result239[92]^and_result239[93]^and_result239[94]^and_result239[95]^and_result239[96]^and_result239[97]^and_result239[98]^and_result239[99]^and_result239[100]^and_result239[101]^and_result239[102]^and_result239[103]^and_result239[104]^and_result239[105]^and_result239[106]^and_result239[107]^and_result239[108]^and_result239[109]^and_result239[110]^and_result239[111]^and_result239[112]^and_result239[113]^and_result239[114]^and_result239[115]^and_result239[116]^and_result239[117]^and_result239[118]^and_result239[119]^and_result239[120]^and_result239[121]^and_result239[122]^and_result239[123]^and_result239[124]^and_result239[125]^and_result239[126]^and_result239[127]^and_result239[128]^and_result239[129]^and_result239[130]^and_result239[131]^and_result239[132]^and_result239[133]^and_result239[134]^and_result239[135]^and_result239[136]^and_result239[137]^and_result239[138]^and_result239[139]^and_result239[140]^and_result239[141]^and_result239[142]^and_result239[143]^and_result239[144]^and_result239[145]^and_result239[146]^and_result239[147]^and_result239[148]^and_result239[149]^and_result239[150]^and_result239[151]^and_result239[152]^and_result239[153]^and_result239[154]^and_result239[155]^and_result239[156]^and_result239[157]^and_result239[158]^and_result239[159]^and_result239[160]^and_result239[161]^and_result239[162]^and_result239[163]^and_result239[164]^and_result239[165]^and_result239[166]^and_result239[167]^and_result239[168]^and_result239[169]^and_result239[170]^and_result239[171]^and_result239[172]^and_result239[173]^and_result239[174]^and_result239[175]^and_result239[176]^and_result239[177]^and_result239[178]^and_result239[179]^and_result239[180]^and_result239[181]^and_result239[182]^and_result239[183]^and_result239[184]^and_result239[185]^and_result239[186]^and_result239[187]^and_result239[188]^and_result239[189]^and_result239[190]^and_result239[191]^and_result239[192]^and_result239[193]^and_result239[194]^and_result239[195]^and_result239[196]^and_result239[197]^and_result239[198]^and_result239[199]^and_result239[200]^and_result239[201]^and_result239[202]^and_result239[203]^and_result239[204]^and_result239[205]^and_result239[206]^and_result239[207]^and_result239[208]^and_result239[209]^and_result239[210]^and_result239[211]^and_result239[212]^and_result239[213]^and_result239[214]^and_result239[215]^and_result239[216]^and_result239[217]^and_result239[218]^and_result239[219]^and_result239[220]^and_result239[221]^and_result239[222]^and_result239[223]^and_result239[224]^and_result239[225]^and_result239[226]^and_result239[227]^and_result239[228]^and_result239[229]^and_result239[230]^and_result239[231]^and_result239[232]^and_result239[233]^and_result239[234]^and_result239[235]^and_result239[236]^and_result239[237]^and_result239[238]^and_result239[239]^and_result239[240]^and_result239[241]^and_result239[242]^and_result239[243]^and_result239[244]^and_result239[245]^and_result239[246]^and_result239[247]^and_result239[248]^and_result239[249]^and_result239[250]^and_result239[251]^and_result239[252]^and_result239[253]^and_result239[254];
assign key[240]=and_result240[0]^and_result240[1]^and_result240[2]^and_result240[3]^and_result240[4]^and_result240[5]^and_result240[6]^and_result240[7]^and_result240[8]^and_result240[9]^and_result240[10]^and_result240[11]^and_result240[12]^and_result240[13]^and_result240[14]^and_result240[15]^and_result240[16]^and_result240[17]^and_result240[18]^and_result240[19]^and_result240[20]^and_result240[21]^and_result240[22]^and_result240[23]^and_result240[24]^and_result240[25]^and_result240[26]^and_result240[27]^and_result240[28]^and_result240[29]^and_result240[30]^and_result240[31]^and_result240[32]^and_result240[33]^and_result240[34]^and_result240[35]^and_result240[36]^and_result240[37]^and_result240[38]^and_result240[39]^and_result240[40]^and_result240[41]^and_result240[42]^and_result240[43]^and_result240[44]^and_result240[45]^and_result240[46]^and_result240[47]^and_result240[48]^and_result240[49]^and_result240[50]^and_result240[51]^and_result240[52]^and_result240[53]^and_result240[54]^and_result240[55]^and_result240[56]^and_result240[57]^and_result240[58]^and_result240[59]^and_result240[60]^and_result240[61]^and_result240[62]^and_result240[63]^and_result240[64]^and_result240[65]^and_result240[66]^and_result240[67]^and_result240[68]^and_result240[69]^and_result240[70]^and_result240[71]^and_result240[72]^and_result240[73]^and_result240[74]^and_result240[75]^and_result240[76]^and_result240[77]^and_result240[78]^and_result240[79]^and_result240[80]^and_result240[81]^and_result240[82]^and_result240[83]^and_result240[84]^and_result240[85]^and_result240[86]^and_result240[87]^and_result240[88]^and_result240[89]^and_result240[90]^and_result240[91]^and_result240[92]^and_result240[93]^and_result240[94]^and_result240[95]^and_result240[96]^and_result240[97]^and_result240[98]^and_result240[99]^and_result240[100]^and_result240[101]^and_result240[102]^and_result240[103]^and_result240[104]^and_result240[105]^and_result240[106]^and_result240[107]^and_result240[108]^and_result240[109]^and_result240[110]^and_result240[111]^and_result240[112]^and_result240[113]^and_result240[114]^and_result240[115]^and_result240[116]^and_result240[117]^and_result240[118]^and_result240[119]^and_result240[120]^and_result240[121]^and_result240[122]^and_result240[123]^and_result240[124]^and_result240[125]^and_result240[126]^and_result240[127]^and_result240[128]^and_result240[129]^and_result240[130]^and_result240[131]^and_result240[132]^and_result240[133]^and_result240[134]^and_result240[135]^and_result240[136]^and_result240[137]^and_result240[138]^and_result240[139]^and_result240[140]^and_result240[141]^and_result240[142]^and_result240[143]^and_result240[144]^and_result240[145]^and_result240[146]^and_result240[147]^and_result240[148]^and_result240[149]^and_result240[150]^and_result240[151]^and_result240[152]^and_result240[153]^and_result240[154]^and_result240[155]^and_result240[156]^and_result240[157]^and_result240[158]^and_result240[159]^and_result240[160]^and_result240[161]^and_result240[162]^and_result240[163]^and_result240[164]^and_result240[165]^and_result240[166]^and_result240[167]^and_result240[168]^and_result240[169]^and_result240[170]^and_result240[171]^and_result240[172]^and_result240[173]^and_result240[174]^and_result240[175]^and_result240[176]^and_result240[177]^and_result240[178]^and_result240[179]^and_result240[180]^and_result240[181]^and_result240[182]^and_result240[183]^and_result240[184]^and_result240[185]^and_result240[186]^and_result240[187]^and_result240[188]^and_result240[189]^and_result240[190]^and_result240[191]^and_result240[192]^and_result240[193]^and_result240[194]^and_result240[195]^and_result240[196]^and_result240[197]^and_result240[198]^and_result240[199]^and_result240[200]^and_result240[201]^and_result240[202]^and_result240[203]^and_result240[204]^and_result240[205]^and_result240[206]^and_result240[207]^and_result240[208]^and_result240[209]^and_result240[210]^and_result240[211]^and_result240[212]^and_result240[213]^and_result240[214]^and_result240[215]^and_result240[216]^and_result240[217]^and_result240[218]^and_result240[219]^and_result240[220]^and_result240[221]^and_result240[222]^and_result240[223]^and_result240[224]^and_result240[225]^and_result240[226]^and_result240[227]^and_result240[228]^and_result240[229]^and_result240[230]^and_result240[231]^and_result240[232]^and_result240[233]^and_result240[234]^and_result240[235]^and_result240[236]^and_result240[237]^and_result240[238]^and_result240[239]^and_result240[240]^and_result240[241]^and_result240[242]^and_result240[243]^and_result240[244]^and_result240[245]^and_result240[246]^and_result240[247]^and_result240[248]^and_result240[249]^and_result240[250]^and_result240[251]^and_result240[252]^and_result240[253]^and_result240[254];
assign key[241]=and_result241[0]^and_result241[1]^and_result241[2]^and_result241[3]^and_result241[4]^and_result241[5]^and_result241[6]^and_result241[7]^and_result241[8]^and_result241[9]^and_result241[10]^and_result241[11]^and_result241[12]^and_result241[13]^and_result241[14]^and_result241[15]^and_result241[16]^and_result241[17]^and_result241[18]^and_result241[19]^and_result241[20]^and_result241[21]^and_result241[22]^and_result241[23]^and_result241[24]^and_result241[25]^and_result241[26]^and_result241[27]^and_result241[28]^and_result241[29]^and_result241[30]^and_result241[31]^and_result241[32]^and_result241[33]^and_result241[34]^and_result241[35]^and_result241[36]^and_result241[37]^and_result241[38]^and_result241[39]^and_result241[40]^and_result241[41]^and_result241[42]^and_result241[43]^and_result241[44]^and_result241[45]^and_result241[46]^and_result241[47]^and_result241[48]^and_result241[49]^and_result241[50]^and_result241[51]^and_result241[52]^and_result241[53]^and_result241[54]^and_result241[55]^and_result241[56]^and_result241[57]^and_result241[58]^and_result241[59]^and_result241[60]^and_result241[61]^and_result241[62]^and_result241[63]^and_result241[64]^and_result241[65]^and_result241[66]^and_result241[67]^and_result241[68]^and_result241[69]^and_result241[70]^and_result241[71]^and_result241[72]^and_result241[73]^and_result241[74]^and_result241[75]^and_result241[76]^and_result241[77]^and_result241[78]^and_result241[79]^and_result241[80]^and_result241[81]^and_result241[82]^and_result241[83]^and_result241[84]^and_result241[85]^and_result241[86]^and_result241[87]^and_result241[88]^and_result241[89]^and_result241[90]^and_result241[91]^and_result241[92]^and_result241[93]^and_result241[94]^and_result241[95]^and_result241[96]^and_result241[97]^and_result241[98]^and_result241[99]^and_result241[100]^and_result241[101]^and_result241[102]^and_result241[103]^and_result241[104]^and_result241[105]^and_result241[106]^and_result241[107]^and_result241[108]^and_result241[109]^and_result241[110]^and_result241[111]^and_result241[112]^and_result241[113]^and_result241[114]^and_result241[115]^and_result241[116]^and_result241[117]^and_result241[118]^and_result241[119]^and_result241[120]^and_result241[121]^and_result241[122]^and_result241[123]^and_result241[124]^and_result241[125]^and_result241[126]^and_result241[127]^and_result241[128]^and_result241[129]^and_result241[130]^and_result241[131]^and_result241[132]^and_result241[133]^and_result241[134]^and_result241[135]^and_result241[136]^and_result241[137]^and_result241[138]^and_result241[139]^and_result241[140]^and_result241[141]^and_result241[142]^and_result241[143]^and_result241[144]^and_result241[145]^and_result241[146]^and_result241[147]^and_result241[148]^and_result241[149]^and_result241[150]^and_result241[151]^and_result241[152]^and_result241[153]^and_result241[154]^and_result241[155]^and_result241[156]^and_result241[157]^and_result241[158]^and_result241[159]^and_result241[160]^and_result241[161]^and_result241[162]^and_result241[163]^and_result241[164]^and_result241[165]^and_result241[166]^and_result241[167]^and_result241[168]^and_result241[169]^and_result241[170]^and_result241[171]^and_result241[172]^and_result241[173]^and_result241[174]^and_result241[175]^and_result241[176]^and_result241[177]^and_result241[178]^and_result241[179]^and_result241[180]^and_result241[181]^and_result241[182]^and_result241[183]^and_result241[184]^and_result241[185]^and_result241[186]^and_result241[187]^and_result241[188]^and_result241[189]^and_result241[190]^and_result241[191]^and_result241[192]^and_result241[193]^and_result241[194]^and_result241[195]^and_result241[196]^and_result241[197]^and_result241[198]^and_result241[199]^and_result241[200]^and_result241[201]^and_result241[202]^and_result241[203]^and_result241[204]^and_result241[205]^and_result241[206]^and_result241[207]^and_result241[208]^and_result241[209]^and_result241[210]^and_result241[211]^and_result241[212]^and_result241[213]^and_result241[214]^and_result241[215]^and_result241[216]^and_result241[217]^and_result241[218]^and_result241[219]^and_result241[220]^and_result241[221]^and_result241[222]^and_result241[223]^and_result241[224]^and_result241[225]^and_result241[226]^and_result241[227]^and_result241[228]^and_result241[229]^and_result241[230]^and_result241[231]^and_result241[232]^and_result241[233]^and_result241[234]^and_result241[235]^and_result241[236]^and_result241[237]^and_result241[238]^and_result241[239]^and_result241[240]^and_result241[241]^and_result241[242]^and_result241[243]^and_result241[244]^and_result241[245]^and_result241[246]^and_result241[247]^and_result241[248]^and_result241[249]^and_result241[250]^and_result241[251]^and_result241[252]^and_result241[253]^and_result241[254];
assign key[242]=and_result242[0]^and_result242[1]^and_result242[2]^and_result242[3]^and_result242[4]^and_result242[5]^and_result242[6]^and_result242[7]^and_result242[8]^and_result242[9]^and_result242[10]^and_result242[11]^and_result242[12]^and_result242[13]^and_result242[14]^and_result242[15]^and_result242[16]^and_result242[17]^and_result242[18]^and_result242[19]^and_result242[20]^and_result242[21]^and_result242[22]^and_result242[23]^and_result242[24]^and_result242[25]^and_result242[26]^and_result242[27]^and_result242[28]^and_result242[29]^and_result242[30]^and_result242[31]^and_result242[32]^and_result242[33]^and_result242[34]^and_result242[35]^and_result242[36]^and_result242[37]^and_result242[38]^and_result242[39]^and_result242[40]^and_result242[41]^and_result242[42]^and_result242[43]^and_result242[44]^and_result242[45]^and_result242[46]^and_result242[47]^and_result242[48]^and_result242[49]^and_result242[50]^and_result242[51]^and_result242[52]^and_result242[53]^and_result242[54]^and_result242[55]^and_result242[56]^and_result242[57]^and_result242[58]^and_result242[59]^and_result242[60]^and_result242[61]^and_result242[62]^and_result242[63]^and_result242[64]^and_result242[65]^and_result242[66]^and_result242[67]^and_result242[68]^and_result242[69]^and_result242[70]^and_result242[71]^and_result242[72]^and_result242[73]^and_result242[74]^and_result242[75]^and_result242[76]^and_result242[77]^and_result242[78]^and_result242[79]^and_result242[80]^and_result242[81]^and_result242[82]^and_result242[83]^and_result242[84]^and_result242[85]^and_result242[86]^and_result242[87]^and_result242[88]^and_result242[89]^and_result242[90]^and_result242[91]^and_result242[92]^and_result242[93]^and_result242[94]^and_result242[95]^and_result242[96]^and_result242[97]^and_result242[98]^and_result242[99]^and_result242[100]^and_result242[101]^and_result242[102]^and_result242[103]^and_result242[104]^and_result242[105]^and_result242[106]^and_result242[107]^and_result242[108]^and_result242[109]^and_result242[110]^and_result242[111]^and_result242[112]^and_result242[113]^and_result242[114]^and_result242[115]^and_result242[116]^and_result242[117]^and_result242[118]^and_result242[119]^and_result242[120]^and_result242[121]^and_result242[122]^and_result242[123]^and_result242[124]^and_result242[125]^and_result242[126]^and_result242[127]^and_result242[128]^and_result242[129]^and_result242[130]^and_result242[131]^and_result242[132]^and_result242[133]^and_result242[134]^and_result242[135]^and_result242[136]^and_result242[137]^and_result242[138]^and_result242[139]^and_result242[140]^and_result242[141]^and_result242[142]^and_result242[143]^and_result242[144]^and_result242[145]^and_result242[146]^and_result242[147]^and_result242[148]^and_result242[149]^and_result242[150]^and_result242[151]^and_result242[152]^and_result242[153]^and_result242[154]^and_result242[155]^and_result242[156]^and_result242[157]^and_result242[158]^and_result242[159]^and_result242[160]^and_result242[161]^and_result242[162]^and_result242[163]^and_result242[164]^and_result242[165]^and_result242[166]^and_result242[167]^and_result242[168]^and_result242[169]^and_result242[170]^and_result242[171]^and_result242[172]^and_result242[173]^and_result242[174]^and_result242[175]^and_result242[176]^and_result242[177]^and_result242[178]^and_result242[179]^and_result242[180]^and_result242[181]^and_result242[182]^and_result242[183]^and_result242[184]^and_result242[185]^and_result242[186]^and_result242[187]^and_result242[188]^and_result242[189]^and_result242[190]^and_result242[191]^and_result242[192]^and_result242[193]^and_result242[194]^and_result242[195]^and_result242[196]^and_result242[197]^and_result242[198]^and_result242[199]^and_result242[200]^and_result242[201]^and_result242[202]^and_result242[203]^and_result242[204]^and_result242[205]^and_result242[206]^and_result242[207]^and_result242[208]^and_result242[209]^and_result242[210]^and_result242[211]^and_result242[212]^and_result242[213]^and_result242[214]^and_result242[215]^and_result242[216]^and_result242[217]^and_result242[218]^and_result242[219]^and_result242[220]^and_result242[221]^and_result242[222]^and_result242[223]^and_result242[224]^and_result242[225]^and_result242[226]^and_result242[227]^and_result242[228]^and_result242[229]^and_result242[230]^and_result242[231]^and_result242[232]^and_result242[233]^and_result242[234]^and_result242[235]^and_result242[236]^and_result242[237]^and_result242[238]^and_result242[239]^and_result242[240]^and_result242[241]^and_result242[242]^and_result242[243]^and_result242[244]^and_result242[245]^and_result242[246]^and_result242[247]^and_result242[248]^and_result242[249]^and_result242[250]^and_result242[251]^and_result242[252]^and_result242[253]^and_result242[254];
assign key[243]=and_result243[0]^and_result243[1]^and_result243[2]^and_result243[3]^and_result243[4]^and_result243[5]^and_result243[6]^and_result243[7]^and_result243[8]^and_result243[9]^and_result243[10]^and_result243[11]^and_result243[12]^and_result243[13]^and_result243[14]^and_result243[15]^and_result243[16]^and_result243[17]^and_result243[18]^and_result243[19]^and_result243[20]^and_result243[21]^and_result243[22]^and_result243[23]^and_result243[24]^and_result243[25]^and_result243[26]^and_result243[27]^and_result243[28]^and_result243[29]^and_result243[30]^and_result243[31]^and_result243[32]^and_result243[33]^and_result243[34]^and_result243[35]^and_result243[36]^and_result243[37]^and_result243[38]^and_result243[39]^and_result243[40]^and_result243[41]^and_result243[42]^and_result243[43]^and_result243[44]^and_result243[45]^and_result243[46]^and_result243[47]^and_result243[48]^and_result243[49]^and_result243[50]^and_result243[51]^and_result243[52]^and_result243[53]^and_result243[54]^and_result243[55]^and_result243[56]^and_result243[57]^and_result243[58]^and_result243[59]^and_result243[60]^and_result243[61]^and_result243[62]^and_result243[63]^and_result243[64]^and_result243[65]^and_result243[66]^and_result243[67]^and_result243[68]^and_result243[69]^and_result243[70]^and_result243[71]^and_result243[72]^and_result243[73]^and_result243[74]^and_result243[75]^and_result243[76]^and_result243[77]^and_result243[78]^and_result243[79]^and_result243[80]^and_result243[81]^and_result243[82]^and_result243[83]^and_result243[84]^and_result243[85]^and_result243[86]^and_result243[87]^and_result243[88]^and_result243[89]^and_result243[90]^and_result243[91]^and_result243[92]^and_result243[93]^and_result243[94]^and_result243[95]^and_result243[96]^and_result243[97]^and_result243[98]^and_result243[99]^and_result243[100]^and_result243[101]^and_result243[102]^and_result243[103]^and_result243[104]^and_result243[105]^and_result243[106]^and_result243[107]^and_result243[108]^and_result243[109]^and_result243[110]^and_result243[111]^and_result243[112]^and_result243[113]^and_result243[114]^and_result243[115]^and_result243[116]^and_result243[117]^and_result243[118]^and_result243[119]^and_result243[120]^and_result243[121]^and_result243[122]^and_result243[123]^and_result243[124]^and_result243[125]^and_result243[126]^and_result243[127]^and_result243[128]^and_result243[129]^and_result243[130]^and_result243[131]^and_result243[132]^and_result243[133]^and_result243[134]^and_result243[135]^and_result243[136]^and_result243[137]^and_result243[138]^and_result243[139]^and_result243[140]^and_result243[141]^and_result243[142]^and_result243[143]^and_result243[144]^and_result243[145]^and_result243[146]^and_result243[147]^and_result243[148]^and_result243[149]^and_result243[150]^and_result243[151]^and_result243[152]^and_result243[153]^and_result243[154]^and_result243[155]^and_result243[156]^and_result243[157]^and_result243[158]^and_result243[159]^and_result243[160]^and_result243[161]^and_result243[162]^and_result243[163]^and_result243[164]^and_result243[165]^and_result243[166]^and_result243[167]^and_result243[168]^and_result243[169]^and_result243[170]^and_result243[171]^and_result243[172]^and_result243[173]^and_result243[174]^and_result243[175]^and_result243[176]^and_result243[177]^and_result243[178]^and_result243[179]^and_result243[180]^and_result243[181]^and_result243[182]^and_result243[183]^and_result243[184]^and_result243[185]^and_result243[186]^and_result243[187]^and_result243[188]^and_result243[189]^and_result243[190]^and_result243[191]^and_result243[192]^and_result243[193]^and_result243[194]^and_result243[195]^and_result243[196]^and_result243[197]^and_result243[198]^and_result243[199]^and_result243[200]^and_result243[201]^and_result243[202]^and_result243[203]^and_result243[204]^and_result243[205]^and_result243[206]^and_result243[207]^and_result243[208]^and_result243[209]^and_result243[210]^and_result243[211]^and_result243[212]^and_result243[213]^and_result243[214]^and_result243[215]^and_result243[216]^and_result243[217]^and_result243[218]^and_result243[219]^and_result243[220]^and_result243[221]^and_result243[222]^and_result243[223]^and_result243[224]^and_result243[225]^and_result243[226]^and_result243[227]^and_result243[228]^and_result243[229]^and_result243[230]^and_result243[231]^and_result243[232]^and_result243[233]^and_result243[234]^and_result243[235]^and_result243[236]^and_result243[237]^and_result243[238]^and_result243[239]^and_result243[240]^and_result243[241]^and_result243[242]^and_result243[243]^and_result243[244]^and_result243[245]^and_result243[246]^and_result243[247]^and_result243[248]^and_result243[249]^and_result243[250]^and_result243[251]^and_result243[252]^and_result243[253]^and_result243[254];
assign key[244]=and_result244[0]^and_result244[1]^and_result244[2]^and_result244[3]^and_result244[4]^and_result244[5]^and_result244[6]^and_result244[7]^and_result244[8]^and_result244[9]^and_result244[10]^and_result244[11]^and_result244[12]^and_result244[13]^and_result244[14]^and_result244[15]^and_result244[16]^and_result244[17]^and_result244[18]^and_result244[19]^and_result244[20]^and_result244[21]^and_result244[22]^and_result244[23]^and_result244[24]^and_result244[25]^and_result244[26]^and_result244[27]^and_result244[28]^and_result244[29]^and_result244[30]^and_result244[31]^and_result244[32]^and_result244[33]^and_result244[34]^and_result244[35]^and_result244[36]^and_result244[37]^and_result244[38]^and_result244[39]^and_result244[40]^and_result244[41]^and_result244[42]^and_result244[43]^and_result244[44]^and_result244[45]^and_result244[46]^and_result244[47]^and_result244[48]^and_result244[49]^and_result244[50]^and_result244[51]^and_result244[52]^and_result244[53]^and_result244[54]^and_result244[55]^and_result244[56]^and_result244[57]^and_result244[58]^and_result244[59]^and_result244[60]^and_result244[61]^and_result244[62]^and_result244[63]^and_result244[64]^and_result244[65]^and_result244[66]^and_result244[67]^and_result244[68]^and_result244[69]^and_result244[70]^and_result244[71]^and_result244[72]^and_result244[73]^and_result244[74]^and_result244[75]^and_result244[76]^and_result244[77]^and_result244[78]^and_result244[79]^and_result244[80]^and_result244[81]^and_result244[82]^and_result244[83]^and_result244[84]^and_result244[85]^and_result244[86]^and_result244[87]^and_result244[88]^and_result244[89]^and_result244[90]^and_result244[91]^and_result244[92]^and_result244[93]^and_result244[94]^and_result244[95]^and_result244[96]^and_result244[97]^and_result244[98]^and_result244[99]^and_result244[100]^and_result244[101]^and_result244[102]^and_result244[103]^and_result244[104]^and_result244[105]^and_result244[106]^and_result244[107]^and_result244[108]^and_result244[109]^and_result244[110]^and_result244[111]^and_result244[112]^and_result244[113]^and_result244[114]^and_result244[115]^and_result244[116]^and_result244[117]^and_result244[118]^and_result244[119]^and_result244[120]^and_result244[121]^and_result244[122]^and_result244[123]^and_result244[124]^and_result244[125]^and_result244[126]^and_result244[127]^and_result244[128]^and_result244[129]^and_result244[130]^and_result244[131]^and_result244[132]^and_result244[133]^and_result244[134]^and_result244[135]^and_result244[136]^and_result244[137]^and_result244[138]^and_result244[139]^and_result244[140]^and_result244[141]^and_result244[142]^and_result244[143]^and_result244[144]^and_result244[145]^and_result244[146]^and_result244[147]^and_result244[148]^and_result244[149]^and_result244[150]^and_result244[151]^and_result244[152]^and_result244[153]^and_result244[154]^and_result244[155]^and_result244[156]^and_result244[157]^and_result244[158]^and_result244[159]^and_result244[160]^and_result244[161]^and_result244[162]^and_result244[163]^and_result244[164]^and_result244[165]^and_result244[166]^and_result244[167]^and_result244[168]^and_result244[169]^and_result244[170]^and_result244[171]^and_result244[172]^and_result244[173]^and_result244[174]^and_result244[175]^and_result244[176]^and_result244[177]^and_result244[178]^and_result244[179]^and_result244[180]^and_result244[181]^and_result244[182]^and_result244[183]^and_result244[184]^and_result244[185]^and_result244[186]^and_result244[187]^and_result244[188]^and_result244[189]^and_result244[190]^and_result244[191]^and_result244[192]^and_result244[193]^and_result244[194]^and_result244[195]^and_result244[196]^and_result244[197]^and_result244[198]^and_result244[199]^and_result244[200]^and_result244[201]^and_result244[202]^and_result244[203]^and_result244[204]^and_result244[205]^and_result244[206]^and_result244[207]^and_result244[208]^and_result244[209]^and_result244[210]^and_result244[211]^and_result244[212]^and_result244[213]^and_result244[214]^and_result244[215]^and_result244[216]^and_result244[217]^and_result244[218]^and_result244[219]^and_result244[220]^and_result244[221]^and_result244[222]^and_result244[223]^and_result244[224]^and_result244[225]^and_result244[226]^and_result244[227]^and_result244[228]^and_result244[229]^and_result244[230]^and_result244[231]^and_result244[232]^and_result244[233]^and_result244[234]^and_result244[235]^and_result244[236]^and_result244[237]^and_result244[238]^and_result244[239]^and_result244[240]^and_result244[241]^and_result244[242]^and_result244[243]^and_result244[244]^and_result244[245]^and_result244[246]^and_result244[247]^and_result244[248]^and_result244[249]^and_result244[250]^and_result244[251]^and_result244[252]^and_result244[253]^and_result244[254];
assign key[245]=and_result245[0]^and_result245[1]^and_result245[2]^and_result245[3]^and_result245[4]^and_result245[5]^and_result245[6]^and_result245[7]^and_result245[8]^and_result245[9]^and_result245[10]^and_result245[11]^and_result245[12]^and_result245[13]^and_result245[14]^and_result245[15]^and_result245[16]^and_result245[17]^and_result245[18]^and_result245[19]^and_result245[20]^and_result245[21]^and_result245[22]^and_result245[23]^and_result245[24]^and_result245[25]^and_result245[26]^and_result245[27]^and_result245[28]^and_result245[29]^and_result245[30]^and_result245[31]^and_result245[32]^and_result245[33]^and_result245[34]^and_result245[35]^and_result245[36]^and_result245[37]^and_result245[38]^and_result245[39]^and_result245[40]^and_result245[41]^and_result245[42]^and_result245[43]^and_result245[44]^and_result245[45]^and_result245[46]^and_result245[47]^and_result245[48]^and_result245[49]^and_result245[50]^and_result245[51]^and_result245[52]^and_result245[53]^and_result245[54]^and_result245[55]^and_result245[56]^and_result245[57]^and_result245[58]^and_result245[59]^and_result245[60]^and_result245[61]^and_result245[62]^and_result245[63]^and_result245[64]^and_result245[65]^and_result245[66]^and_result245[67]^and_result245[68]^and_result245[69]^and_result245[70]^and_result245[71]^and_result245[72]^and_result245[73]^and_result245[74]^and_result245[75]^and_result245[76]^and_result245[77]^and_result245[78]^and_result245[79]^and_result245[80]^and_result245[81]^and_result245[82]^and_result245[83]^and_result245[84]^and_result245[85]^and_result245[86]^and_result245[87]^and_result245[88]^and_result245[89]^and_result245[90]^and_result245[91]^and_result245[92]^and_result245[93]^and_result245[94]^and_result245[95]^and_result245[96]^and_result245[97]^and_result245[98]^and_result245[99]^and_result245[100]^and_result245[101]^and_result245[102]^and_result245[103]^and_result245[104]^and_result245[105]^and_result245[106]^and_result245[107]^and_result245[108]^and_result245[109]^and_result245[110]^and_result245[111]^and_result245[112]^and_result245[113]^and_result245[114]^and_result245[115]^and_result245[116]^and_result245[117]^and_result245[118]^and_result245[119]^and_result245[120]^and_result245[121]^and_result245[122]^and_result245[123]^and_result245[124]^and_result245[125]^and_result245[126]^and_result245[127]^and_result245[128]^and_result245[129]^and_result245[130]^and_result245[131]^and_result245[132]^and_result245[133]^and_result245[134]^and_result245[135]^and_result245[136]^and_result245[137]^and_result245[138]^and_result245[139]^and_result245[140]^and_result245[141]^and_result245[142]^and_result245[143]^and_result245[144]^and_result245[145]^and_result245[146]^and_result245[147]^and_result245[148]^and_result245[149]^and_result245[150]^and_result245[151]^and_result245[152]^and_result245[153]^and_result245[154]^and_result245[155]^and_result245[156]^and_result245[157]^and_result245[158]^and_result245[159]^and_result245[160]^and_result245[161]^and_result245[162]^and_result245[163]^and_result245[164]^and_result245[165]^and_result245[166]^and_result245[167]^and_result245[168]^and_result245[169]^and_result245[170]^and_result245[171]^and_result245[172]^and_result245[173]^and_result245[174]^and_result245[175]^and_result245[176]^and_result245[177]^and_result245[178]^and_result245[179]^and_result245[180]^and_result245[181]^and_result245[182]^and_result245[183]^and_result245[184]^and_result245[185]^and_result245[186]^and_result245[187]^and_result245[188]^and_result245[189]^and_result245[190]^and_result245[191]^and_result245[192]^and_result245[193]^and_result245[194]^and_result245[195]^and_result245[196]^and_result245[197]^and_result245[198]^and_result245[199]^and_result245[200]^and_result245[201]^and_result245[202]^and_result245[203]^and_result245[204]^and_result245[205]^and_result245[206]^and_result245[207]^and_result245[208]^and_result245[209]^and_result245[210]^and_result245[211]^and_result245[212]^and_result245[213]^and_result245[214]^and_result245[215]^and_result245[216]^and_result245[217]^and_result245[218]^and_result245[219]^and_result245[220]^and_result245[221]^and_result245[222]^and_result245[223]^and_result245[224]^and_result245[225]^and_result245[226]^and_result245[227]^and_result245[228]^and_result245[229]^and_result245[230]^and_result245[231]^and_result245[232]^and_result245[233]^and_result245[234]^and_result245[235]^and_result245[236]^and_result245[237]^and_result245[238]^and_result245[239]^and_result245[240]^and_result245[241]^and_result245[242]^and_result245[243]^and_result245[244]^and_result245[245]^and_result245[246]^and_result245[247]^and_result245[248]^and_result245[249]^and_result245[250]^and_result245[251]^and_result245[252]^and_result245[253]^and_result245[254];
assign key[246]=and_result246[0]^and_result246[1]^and_result246[2]^and_result246[3]^and_result246[4]^and_result246[5]^and_result246[6]^and_result246[7]^and_result246[8]^and_result246[9]^and_result246[10]^and_result246[11]^and_result246[12]^and_result246[13]^and_result246[14]^and_result246[15]^and_result246[16]^and_result246[17]^and_result246[18]^and_result246[19]^and_result246[20]^and_result246[21]^and_result246[22]^and_result246[23]^and_result246[24]^and_result246[25]^and_result246[26]^and_result246[27]^and_result246[28]^and_result246[29]^and_result246[30]^and_result246[31]^and_result246[32]^and_result246[33]^and_result246[34]^and_result246[35]^and_result246[36]^and_result246[37]^and_result246[38]^and_result246[39]^and_result246[40]^and_result246[41]^and_result246[42]^and_result246[43]^and_result246[44]^and_result246[45]^and_result246[46]^and_result246[47]^and_result246[48]^and_result246[49]^and_result246[50]^and_result246[51]^and_result246[52]^and_result246[53]^and_result246[54]^and_result246[55]^and_result246[56]^and_result246[57]^and_result246[58]^and_result246[59]^and_result246[60]^and_result246[61]^and_result246[62]^and_result246[63]^and_result246[64]^and_result246[65]^and_result246[66]^and_result246[67]^and_result246[68]^and_result246[69]^and_result246[70]^and_result246[71]^and_result246[72]^and_result246[73]^and_result246[74]^and_result246[75]^and_result246[76]^and_result246[77]^and_result246[78]^and_result246[79]^and_result246[80]^and_result246[81]^and_result246[82]^and_result246[83]^and_result246[84]^and_result246[85]^and_result246[86]^and_result246[87]^and_result246[88]^and_result246[89]^and_result246[90]^and_result246[91]^and_result246[92]^and_result246[93]^and_result246[94]^and_result246[95]^and_result246[96]^and_result246[97]^and_result246[98]^and_result246[99]^and_result246[100]^and_result246[101]^and_result246[102]^and_result246[103]^and_result246[104]^and_result246[105]^and_result246[106]^and_result246[107]^and_result246[108]^and_result246[109]^and_result246[110]^and_result246[111]^and_result246[112]^and_result246[113]^and_result246[114]^and_result246[115]^and_result246[116]^and_result246[117]^and_result246[118]^and_result246[119]^and_result246[120]^and_result246[121]^and_result246[122]^and_result246[123]^and_result246[124]^and_result246[125]^and_result246[126]^and_result246[127]^and_result246[128]^and_result246[129]^and_result246[130]^and_result246[131]^and_result246[132]^and_result246[133]^and_result246[134]^and_result246[135]^and_result246[136]^and_result246[137]^and_result246[138]^and_result246[139]^and_result246[140]^and_result246[141]^and_result246[142]^and_result246[143]^and_result246[144]^and_result246[145]^and_result246[146]^and_result246[147]^and_result246[148]^and_result246[149]^and_result246[150]^and_result246[151]^and_result246[152]^and_result246[153]^and_result246[154]^and_result246[155]^and_result246[156]^and_result246[157]^and_result246[158]^and_result246[159]^and_result246[160]^and_result246[161]^and_result246[162]^and_result246[163]^and_result246[164]^and_result246[165]^and_result246[166]^and_result246[167]^and_result246[168]^and_result246[169]^and_result246[170]^and_result246[171]^and_result246[172]^and_result246[173]^and_result246[174]^and_result246[175]^and_result246[176]^and_result246[177]^and_result246[178]^and_result246[179]^and_result246[180]^and_result246[181]^and_result246[182]^and_result246[183]^and_result246[184]^and_result246[185]^and_result246[186]^and_result246[187]^and_result246[188]^and_result246[189]^and_result246[190]^and_result246[191]^and_result246[192]^and_result246[193]^and_result246[194]^and_result246[195]^and_result246[196]^and_result246[197]^and_result246[198]^and_result246[199]^and_result246[200]^and_result246[201]^and_result246[202]^and_result246[203]^and_result246[204]^and_result246[205]^and_result246[206]^and_result246[207]^and_result246[208]^and_result246[209]^and_result246[210]^and_result246[211]^and_result246[212]^and_result246[213]^and_result246[214]^and_result246[215]^and_result246[216]^and_result246[217]^and_result246[218]^and_result246[219]^and_result246[220]^and_result246[221]^and_result246[222]^and_result246[223]^and_result246[224]^and_result246[225]^and_result246[226]^and_result246[227]^and_result246[228]^and_result246[229]^and_result246[230]^and_result246[231]^and_result246[232]^and_result246[233]^and_result246[234]^and_result246[235]^and_result246[236]^and_result246[237]^and_result246[238]^and_result246[239]^and_result246[240]^and_result246[241]^and_result246[242]^and_result246[243]^and_result246[244]^and_result246[245]^and_result246[246]^and_result246[247]^and_result246[248]^and_result246[249]^and_result246[250]^and_result246[251]^and_result246[252]^and_result246[253]^and_result246[254];
assign key[247]=and_result247[0]^and_result247[1]^and_result247[2]^and_result247[3]^and_result247[4]^and_result247[5]^and_result247[6]^and_result247[7]^and_result247[8]^and_result247[9]^and_result247[10]^and_result247[11]^and_result247[12]^and_result247[13]^and_result247[14]^and_result247[15]^and_result247[16]^and_result247[17]^and_result247[18]^and_result247[19]^and_result247[20]^and_result247[21]^and_result247[22]^and_result247[23]^and_result247[24]^and_result247[25]^and_result247[26]^and_result247[27]^and_result247[28]^and_result247[29]^and_result247[30]^and_result247[31]^and_result247[32]^and_result247[33]^and_result247[34]^and_result247[35]^and_result247[36]^and_result247[37]^and_result247[38]^and_result247[39]^and_result247[40]^and_result247[41]^and_result247[42]^and_result247[43]^and_result247[44]^and_result247[45]^and_result247[46]^and_result247[47]^and_result247[48]^and_result247[49]^and_result247[50]^and_result247[51]^and_result247[52]^and_result247[53]^and_result247[54]^and_result247[55]^and_result247[56]^and_result247[57]^and_result247[58]^and_result247[59]^and_result247[60]^and_result247[61]^and_result247[62]^and_result247[63]^and_result247[64]^and_result247[65]^and_result247[66]^and_result247[67]^and_result247[68]^and_result247[69]^and_result247[70]^and_result247[71]^and_result247[72]^and_result247[73]^and_result247[74]^and_result247[75]^and_result247[76]^and_result247[77]^and_result247[78]^and_result247[79]^and_result247[80]^and_result247[81]^and_result247[82]^and_result247[83]^and_result247[84]^and_result247[85]^and_result247[86]^and_result247[87]^and_result247[88]^and_result247[89]^and_result247[90]^and_result247[91]^and_result247[92]^and_result247[93]^and_result247[94]^and_result247[95]^and_result247[96]^and_result247[97]^and_result247[98]^and_result247[99]^and_result247[100]^and_result247[101]^and_result247[102]^and_result247[103]^and_result247[104]^and_result247[105]^and_result247[106]^and_result247[107]^and_result247[108]^and_result247[109]^and_result247[110]^and_result247[111]^and_result247[112]^and_result247[113]^and_result247[114]^and_result247[115]^and_result247[116]^and_result247[117]^and_result247[118]^and_result247[119]^and_result247[120]^and_result247[121]^and_result247[122]^and_result247[123]^and_result247[124]^and_result247[125]^and_result247[126]^and_result247[127]^and_result247[128]^and_result247[129]^and_result247[130]^and_result247[131]^and_result247[132]^and_result247[133]^and_result247[134]^and_result247[135]^and_result247[136]^and_result247[137]^and_result247[138]^and_result247[139]^and_result247[140]^and_result247[141]^and_result247[142]^and_result247[143]^and_result247[144]^and_result247[145]^and_result247[146]^and_result247[147]^and_result247[148]^and_result247[149]^and_result247[150]^and_result247[151]^and_result247[152]^and_result247[153]^and_result247[154]^and_result247[155]^and_result247[156]^and_result247[157]^and_result247[158]^and_result247[159]^and_result247[160]^and_result247[161]^and_result247[162]^and_result247[163]^and_result247[164]^and_result247[165]^and_result247[166]^and_result247[167]^and_result247[168]^and_result247[169]^and_result247[170]^and_result247[171]^and_result247[172]^and_result247[173]^and_result247[174]^and_result247[175]^and_result247[176]^and_result247[177]^and_result247[178]^and_result247[179]^and_result247[180]^and_result247[181]^and_result247[182]^and_result247[183]^and_result247[184]^and_result247[185]^and_result247[186]^and_result247[187]^and_result247[188]^and_result247[189]^and_result247[190]^and_result247[191]^and_result247[192]^and_result247[193]^and_result247[194]^and_result247[195]^and_result247[196]^and_result247[197]^and_result247[198]^and_result247[199]^and_result247[200]^and_result247[201]^and_result247[202]^and_result247[203]^and_result247[204]^and_result247[205]^and_result247[206]^and_result247[207]^and_result247[208]^and_result247[209]^and_result247[210]^and_result247[211]^and_result247[212]^and_result247[213]^and_result247[214]^and_result247[215]^and_result247[216]^and_result247[217]^and_result247[218]^and_result247[219]^and_result247[220]^and_result247[221]^and_result247[222]^and_result247[223]^and_result247[224]^and_result247[225]^and_result247[226]^and_result247[227]^and_result247[228]^and_result247[229]^and_result247[230]^and_result247[231]^and_result247[232]^and_result247[233]^and_result247[234]^and_result247[235]^and_result247[236]^and_result247[237]^and_result247[238]^and_result247[239]^and_result247[240]^and_result247[241]^and_result247[242]^and_result247[243]^and_result247[244]^and_result247[245]^and_result247[246]^and_result247[247]^and_result247[248]^and_result247[249]^and_result247[250]^and_result247[251]^and_result247[252]^and_result247[253]^and_result247[254];
assign key[248]=and_result248[0]^and_result248[1]^and_result248[2]^and_result248[3]^and_result248[4]^and_result248[5]^and_result248[6]^and_result248[7]^and_result248[8]^and_result248[9]^and_result248[10]^and_result248[11]^and_result248[12]^and_result248[13]^and_result248[14]^and_result248[15]^and_result248[16]^and_result248[17]^and_result248[18]^and_result248[19]^and_result248[20]^and_result248[21]^and_result248[22]^and_result248[23]^and_result248[24]^and_result248[25]^and_result248[26]^and_result248[27]^and_result248[28]^and_result248[29]^and_result248[30]^and_result248[31]^and_result248[32]^and_result248[33]^and_result248[34]^and_result248[35]^and_result248[36]^and_result248[37]^and_result248[38]^and_result248[39]^and_result248[40]^and_result248[41]^and_result248[42]^and_result248[43]^and_result248[44]^and_result248[45]^and_result248[46]^and_result248[47]^and_result248[48]^and_result248[49]^and_result248[50]^and_result248[51]^and_result248[52]^and_result248[53]^and_result248[54]^and_result248[55]^and_result248[56]^and_result248[57]^and_result248[58]^and_result248[59]^and_result248[60]^and_result248[61]^and_result248[62]^and_result248[63]^and_result248[64]^and_result248[65]^and_result248[66]^and_result248[67]^and_result248[68]^and_result248[69]^and_result248[70]^and_result248[71]^and_result248[72]^and_result248[73]^and_result248[74]^and_result248[75]^and_result248[76]^and_result248[77]^and_result248[78]^and_result248[79]^and_result248[80]^and_result248[81]^and_result248[82]^and_result248[83]^and_result248[84]^and_result248[85]^and_result248[86]^and_result248[87]^and_result248[88]^and_result248[89]^and_result248[90]^and_result248[91]^and_result248[92]^and_result248[93]^and_result248[94]^and_result248[95]^and_result248[96]^and_result248[97]^and_result248[98]^and_result248[99]^and_result248[100]^and_result248[101]^and_result248[102]^and_result248[103]^and_result248[104]^and_result248[105]^and_result248[106]^and_result248[107]^and_result248[108]^and_result248[109]^and_result248[110]^and_result248[111]^and_result248[112]^and_result248[113]^and_result248[114]^and_result248[115]^and_result248[116]^and_result248[117]^and_result248[118]^and_result248[119]^and_result248[120]^and_result248[121]^and_result248[122]^and_result248[123]^and_result248[124]^and_result248[125]^and_result248[126]^and_result248[127]^and_result248[128]^and_result248[129]^and_result248[130]^and_result248[131]^and_result248[132]^and_result248[133]^and_result248[134]^and_result248[135]^and_result248[136]^and_result248[137]^and_result248[138]^and_result248[139]^and_result248[140]^and_result248[141]^and_result248[142]^and_result248[143]^and_result248[144]^and_result248[145]^and_result248[146]^and_result248[147]^and_result248[148]^and_result248[149]^and_result248[150]^and_result248[151]^and_result248[152]^and_result248[153]^and_result248[154]^and_result248[155]^and_result248[156]^and_result248[157]^and_result248[158]^and_result248[159]^and_result248[160]^and_result248[161]^and_result248[162]^and_result248[163]^and_result248[164]^and_result248[165]^and_result248[166]^and_result248[167]^and_result248[168]^and_result248[169]^and_result248[170]^and_result248[171]^and_result248[172]^and_result248[173]^and_result248[174]^and_result248[175]^and_result248[176]^and_result248[177]^and_result248[178]^and_result248[179]^and_result248[180]^and_result248[181]^and_result248[182]^and_result248[183]^and_result248[184]^and_result248[185]^and_result248[186]^and_result248[187]^and_result248[188]^and_result248[189]^and_result248[190]^and_result248[191]^and_result248[192]^and_result248[193]^and_result248[194]^and_result248[195]^and_result248[196]^and_result248[197]^and_result248[198]^and_result248[199]^and_result248[200]^and_result248[201]^and_result248[202]^and_result248[203]^and_result248[204]^and_result248[205]^and_result248[206]^and_result248[207]^and_result248[208]^and_result248[209]^and_result248[210]^and_result248[211]^and_result248[212]^and_result248[213]^and_result248[214]^and_result248[215]^and_result248[216]^and_result248[217]^and_result248[218]^and_result248[219]^and_result248[220]^and_result248[221]^and_result248[222]^and_result248[223]^and_result248[224]^and_result248[225]^and_result248[226]^and_result248[227]^and_result248[228]^and_result248[229]^and_result248[230]^and_result248[231]^and_result248[232]^and_result248[233]^and_result248[234]^and_result248[235]^and_result248[236]^and_result248[237]^and_result248[238]^and_result248[239]^and_result248[240]^and_result248[241]^and_result248[242]^and_result248[243]^and_result248[244]^and_result248[245]^and_result248[246]^and_result248[247]^and_result248[248]^and_result248[249]^and_result248[250]^and_result248[251]^and_result248[252]^and_result248[253]^and_result248[254];
assign key[249]=and_result249[0]^and_result249[1]^and_result249[2]^and_result249[3]^and_result249[4]^and_result249[5]^and_result249[6]^and_result249[7]^and_result249[8]^and_result249[9]^and_result249[10]^and_result249[11]^and_result249[12]^and_result249[13]^and_result249[14]^and_result249[15]^and_result249[16]^and_result249[17]^and_result249[18]^and_result249[19]^and_result249[20]^and_result249[21]^and_result249[22]^and_result249[23]^and_result249[24]^and_result249[25]^and_result249[26]^and_result249[27]^and_result249[28]^and_result249[29]^and_result249[30]^and_result249[31]^and_result249[32]^and_result249[33]^and_result249[34]^and_result249[35]^and_result249[36]^and_result249[37]^and_result249[38]^and_result249[39]^and_result249[40]^and_result249[41]^and_result249[42]^and_result249[43]^and_result249[44]^and_result249[45]^and_result249[46]^and_result249[47]^and_result249[48]^and_result249[49]^and_result249[50]^and_result249[51]^and_result249[52]^and_result249[53]^and_result249[54]^and_result249[55]^and_result249[56]^and_result249[57]^and_result249[58]^and_result249[59]^and_result249[60]^and_result249[61]^and_result249[62]^and_result249[63]^and_result249[64]^and_result249[65]^and_result249[66]^and_result249[67]^and_result249[68]^and_result249[69]^and_result249[70]^and_result249[71]^and_result249[72]^and_result249[73]^and_result249[74]^and_result249[75]^and_result249[76]^and_result249[77]^and_result249[78]^and_result249[79]^and_result249[80]^and_result249[81]^and_result249[82]^and_result249[83]^and_result249[84]^and_result249[85]^and_result249[86]^and_result249[87]^and_result249[88]^and_result249[89]^and_result249[90]^and_result249[91]^and_result249[92]^and_result249[93]^and_result249[94]^and_result249[95]^and_result249[96]^and_result249[97]^and_result249[98]^and_result249[99]^and_result249[100]^and_result249[101]^and_result249[102]^and_result249[103]^and_result249[104]^and_result249[105]^and_result249[106]^and_result249[107]^and_result249[108]^and_result249[109]^and_result249[110]^and_result249[111]^and_result249[112]^and_result249[113]^and_result249[114]^and_result249[115]^and_result249[116]^and_result249[117]^and_result249[118]^and_result249[119]^and_result249[120]^and_result249[121]^and_result249[122]^and_result249[123]^and_result249[124]^and_result249[125]^and_result249[126]^and_result249[127]^and_result249[128]^and_result249[129]^and_result249[130]^and_result249[131]^and_result249[132]^and_result249[133]^and_result249[134]^and_result249[135]^and_result249[136]^and_result249[137]^and_result249[138]^and_result249[139]^and_result249[140]^and_result249[141]^and_result249[142]^and_result249[143]^and_result249[144]^and_result249[145]^and_result249[146]^and_result249[147]^and_result249[148]^and_result249[149]^and_result249[150]^and_result249[151]^and_result249[152]^and_result249[153]^and_result249[154]^and_result249[155]^and_result249[156]^and_result249[157]^and_result249[158]^and_result249[159]^and_result249[160]^and_result249[161]^and_result249[162]^and_result249[163]^and_result249[164]^and_result249[165]^and_result249[166]^and_result249[167]^and_result249[168]^and_result249[169]^and_result249[170]^and_result249[171]^and_result249[172]^and_result249[173]^and_result249[174]^and_result249[175]^and_result249[176]^and_result249[177]^and_result249[178]^and_result249[179]^and_result249[180]^and_result249[181]^and_result249[182]^and_result249[183]^and_result249[184]^and_result249[185]^and_result249[186]^and_result249[187]^and_result249[188]^and_result249[189]^and_result249[190]^and_result249[191]^and_result249[192]^and_result249[193]^and_result249[194]^and_result249[195]^and_result249[196]^and_result249[197]^and_result249[198]^and_result249[199]^and_result249[200]^and_result249[201]^and_result249[202]^and_result249[203]^and_result249[204]^and_result249[205]^and_result249[206]^and_result249[207]^and_result249[208]^and_result249[209]^and_result249[210]^and_result249[211]^and_result249[212]^and_result249[213]^and_result249[214]^and_result249[215]^and_result249[216]^and_result249[217]^and_result249[218]^and_result249[219]^and_result249[220]^and_result249[221]^and_result249[222]^and_result249[223]^and_result249[224]^and_result249[225]^and_result249[226]^and_result249[227]^and_result249[228]^and_result249[229]^and_result249[230]^and_result249[231]^and_result249[232]^and_result249[233]^and_result249[234]^and_result249[235]^and_result249[236]^and_result249[237]^and_result249[238]^and_result249[239]^and_result249[240]^and_result249[241]^and_result249[242]^and_result249[243]^and_result249[244]^and_result249[245]^and_result249[246]^and_result249[247]^and_result249[248]^and_result249[249]^and_result249[250]^and_result249[251]^and_result249[252]^and_result249[253]^and_result249[254];
assign key[250]=and_result250[0]^and_result250[1]^and_result250[2]^and_result250[3]^and_result250[4]^and_result250[5]^and_result250[6]^and_result250[7]^and_result250[8]^and_result250[9]^and_result250[10]^and_result250[11]^and_result250[12]^and_result250[13]^and_result250[14]^and_result250[15]^and_result250[16]^and_result250[17]^and_result250[18]^and_result250[19]^and_result250[20]^and_result250[21]^and_result250[22]^and_result250[23]^and_result250[24]^and_result250[25]^and_result250[26]^and_result250[27]^and_result250[28]^and_result250[29]^and_result250[30]^and_result250[31]^and_result250[32]^and_result250[33]^and_result250[34]^and_result250[35]^and_result250[36]^and_result250[37]^and_result250[38]^and_result250[39]^and_result250[40]^and_result250[41]^and_result250[42]^and_result250[43]^and_result250[44]^and_result250[45]^and_result250[46]^and_result250[47]^and_result250[48]^and_result250[49]^and_result250[50]^and_result250[51]^and_result250[52]^and_result250[53]^and_result250[54]^and_result250[55]^and_result250[56]^and_result250[57]^and_result250[58]^and_result250[59]^and_result250[60]^and_result250[61]^and_result250[62]^and_result250[63]^and_result250[64]^and_result250[65]^and_result250[66]^and_result250[67]^and_result250[68]^and_result250[69]^and_result250[70]^and_result250[71]^and_result250[72]^and_result250[73]^and_result250[74]^and_result250[75]^and_result250[76]^and_result250[77]^and_result250[78]^and_result250[79]^and_result250[80]^and_result250[81]^and_result250[82]^and_result250[83]^and_result250[84]^and_result250[85]^and_result250[86]^and_result250[87]^and_result250[88]^and_result250[89]^and_result250[90]^and_result250[91]^and_result250[92]^and_result250[93]^and_result250[94]^and_result250[95]^and_result250[96]^and_result250[97]^and_result250[98]^and_result250[99]^and_result250[100]^and_result250[101]^and_result250[102]^and_result250[103]^and_result250[104]^and_result250[105]^and_result250[106]^and_result250[107]^and_result250[108]^and_result250[109]^and_result250[110]^and_result250[111]^and_result250[112]^and_result250[113]^and_result250[114]^and_result250[115]^and_result250[116]^and_result250[117]^and_result250[118]^and_result250[119]^and_result250[120]^and_result250[121]^and_result250[122]^and_result250[123]^and_result250[124]^and_result250[125]^and_result250[126]^and_result250[127]^and_result250[128]^and_result250[129]^and_result250[130]^and_result250[131]^and_result250[132]^and_result250[133]^and_result250[134]^and_result250[135]^and_result250[136]^and_result250[137]^and_result250[138]^and_result250[139]^and_result250[140]^and_result250[141]^and_result250[142]^and_result250[143]^and_result250[144]^and_result250[145]^and_result250[146]^and_result250[147]^and_result250[148]^and_result250[149]^and_result250[150]^and_result250[151]^and_result250[152]^and_result250[153]^and_result250[154]^and_result250[155]^and_result250[156]^and_result250[157]^and_result250[158]^and_result250[159]^and_result250[160]^and_result250[161]^and_result250[162]^and_result250[163]^and_result250[164]^and_result250[165]^and_result250[166]^and_result250[167]^and_result250[168]^and_result250[169]^and_result250[170]^and_result250[171]^and_result250[172]^and_result250[173]^and_result250[174]^and_result250[175]^and_result250[176]^and_result250[177]^and_result250[178]^and_result250[179]^and_result250[180]^and_result250[181]^and_result250[182]^and_result250[183]^and_result250[184]^and_result250[185]^and_result250[186]^and_result250[187]^and_result250[188]^and_result250[189]^and_result250[190]^and_result250[191]^and_result250[192]^and_result250[193]^and_result250[194]^and_result250[195]^and_result250[196]^and_result250[197]^and_result250[198]^and_result250[199]^and_result250[200]^and_result250[201]^and_result250[202]^and_result250[203]^and_result250[204]^and_result250[205]^and_result250[206]^and_result250[207]^and_result250[208]^and_result250[209]^and_result250[210]^and_result250[211]^and_result250[212]^and_result250[213]^and_result250[214]^and_result250[215]^and_result250[216]^and_result250[217]^and_result250[218]^and_result250[219]^and_result250[220]^and_result250[221]^and_result250[222]^and_result250[223]^and_result250[224]^and_result250[225]^and_result250[226]^and_result250[227]^and_result250[228]^and_result250[229]^and_result250[230]^and_result250[231]^and_result250[232]^and_result250[233]^and_result250[234]^and_result250[235]^and_result250[236]^and_result250[237]^and_result250[238]^and_result250[239]^and_result250[240]^and_result250[241]^and_result250[242]^and_result250[243]^and_result250[244]^and_result250[245]^and_result250[246]^and_result250[247]^and_result250[248]^and_result250[249]^and_result250[250]^and_result250[251]^and_result250[252]^and_result250[253]^and_result250[254];
assign key[251]=and_result251[0]^and_result251[1]^and_result251[2]^and_result251[3]^and_result251[4]^and_result251[5]^and_result251[6]^and_result251[7]^and_result251[8]^and_result251[9]^and_result251[10]^and_result251[11]^and_result251[12]^and_result251[13]^and_result251[14]^and_result251[15]^and_result251[16]^and_result251[17]^and_result251[18]^and_result251[19]^and_result251[20]^and_result251[21]^and_result251[22]^and_result251[23]^and_result251[24]^and_result251[25]^and_result251[26]^and_result251[27]^and_result251[28]^and_result251[29]^and_result251[30]^and_result251[31]^and_result251[32]^and_result251[33]^and_result251[34]^and_result251[35]^and_result251[36]^and_result251[37]^and_result251[38]^and_result251[39]^and_result251[40]^and_result251[41]^and_result251[42]^and_result251[43]^and_result251[44]^and_result251[45]^and_result251[46]^and_result251[47]^and_result251[48]^and_result251[49]^and_result251[50]^and_result251[51]^and_result251[52]^and_result251[53]^and_result251[54]^and_result251[55]^and_result251[56]^and_result251[57]^and_result251[58]^and_result251[59]^and_result251[60]^and_result251[61]^and_result251[62]^and_result251[63]^and_result251[64]^and_result251[65]^and_result251[66]^and_result251[67]^and_result251[68]^and_result251[69]^and_result251[70]^and_result251[71]^and_result251[72]^and_result251[73]^and_result251[74]^and_result251[75]^and_result251[76]^and_result251[77]^and_result251[78]^and_result251[79]^and_result251[80]^and_result251[81]^and_result251[82]^and_result251[83]^and_result251[84]^and_result251[85]^and_result251[86]^and_result251[87]^and_result251[88]^and_result251[89]^and_result251[90]^and_result251[91]^and_result251[92]^and_result251[93]^and_result251[94]^and_result251[95]^and_result251[96]^and_result251[97]^and_result251[98]^and_result251[99]^and_result251[100]^and_result251[101]^and_result251[102]^and_result251[103]^and_result251[104]^and_result251[105]^and_result251[106]^and_result251[107]^and_result251[108]^and_result251[109]^and_result251[110]^and_result251[111]^and_result251[112]^and_result251[113]^and_result251[114]^and_result251[115]^and_result251[116]^and_result251[117]^and_result251[118]^and_result251[119]^and_result251[120]^and_result251[121]^and_result251[122]^and_result251[123]^and_result251[124]^and_result251[125]^and_result251[126]^and_result251[127]^and_result251[128]^and_result251[129]^and_result251[130]^and_result251[131]^and_result251[132]^and_result251[133]^and_result251[134]^and_result251[135]^and_result251[136]^and_result251[137]^and_result251[138]^and_result251[139]^and_result251[140]^and_result251[141]^and_result251[142]^and_result251[143]^and_result251[144]^and_result251[145]^and_result251[146]^and_result251[147]^and_result251[148]^and_result251[149]^and_result251[150]^and_result251[151]^and_result251[152]^and_result251[153]^and_result251[154]^and_result251[155]^and_result251[156]^and_result251[157]^and_result251[158]^and_result251[159]^and_result251[160]^and_result251[161]^and_result251[162]^and_result251[163]^and_result251[164]^and_result251[165]^and_result251[166]^and_result251[167]^and_result251[168]^and_result251[169]^and_result251[170]^and_result251[171]^and_result251[172]^and_result251[173]^and_result251[174]^and_result251[175]^and_result251[176]^and_result251[177]^and_result251[178]^and_result251[179]^and_result251[180]^and_result251[181]^and_result251[182]^and_result251[183]^and_result251[184]^and_result251[185]^and_result251[186]^and_result251[187]^and_result251[188]^and_result251[189]^and_result251[190]^and_result251[191]^and_result251[192]^and_result251[193]^and_result251[194]^and_result251[195]^and_result251[196]^and_result251[197]^and_result251[198]^and_result251[199]^and_result251[200]^and_result251[201]^and_result251[202]^and_result251[203]^and_result251[204]^and_result251[205]^and_result251[206]^and_result251[207]^and_result251[208]^and_result251[209]^and_result251[210]^and_result251[211]^and_result251[212]^and_result251[213]^and_result251[214]^and_result251[215]^and_result251[216]^and_result251[217]^and_result251[218]^and_result251[219]^and_result251[220]^and_result251[221]^and_result251[222]^and_result251[223]^and_result251[224]^and_result251[225]^and_result251[226]^and_result251[227]^and_result251[228]^and_result251[229]^and_result251[230]^and_result251[231]^and_result251[232]^and_result251[233]^and_result251[234]^and_result251[235]^and_result251[236]^and_result251[237]^and_result251[238]^and_result251[239]^and_result251[240]^and_result251[241]^and_result251[242]^and_result251[243]^and_result251[244]^and_result251[245]^and_result251[246]^and_result251[247]^and_result251[248]^and_result251[249]^and_result251[250]^and_result251[251]^and_result251[252]^and_result251[253]^and_result251[254];
assign key[252]=and_result252[0]^and_result252[1]^and_result252[2]^and_result252[3]^and_result252[4]^and_result252[5]^and_result252[6]^and_result252[7]^and_result252[8]^and_result252[9]^and_result252[10]^and_result252[11]^and_result252[12]^and_result252[13]^and_result252[14]^and_result252[15]^and_result252[16]^and_result252[17]^and_result252[18]^and_result252[19]^and_result252[20]^and_result252[21]^and_result252[22]^and_result252[23]^and_result252[24]^and_result252[25]^and_result252[26]^and_result252[27]^and_result252[28]^and_result252[29]^and_result252[30]^and_result252[31]^and_result252[32]^and_result252[33]^and_result252[34]^and_result252[35]^and_result252[36]^and_result252[37]^and_result252[38]^and_result252[39]^and_result252[40]^and_result252[41]^and_result252[42]^and_result252[43]^and_result252[44]^and_result252[45]^and_result252[46]^and_result252[47]^and_result252[48]^and_result252[49]^and_result252[50]^and_result252[51]^and_result252[52]^and_result252[53]^and_result252[54]^and_result252[55]^and_result252[56]^and_result252[57]^and_result252[58]^and_result252[59]^and_result252[60]^and_result252[61]^and_result252[62]^and_result252[63]^and_result252[64]^and_result252[65]^and_result252[66]^and_result252[67]^and_result252[68]^and_result252[69]^and_result252[70]^and_result252[71]^and_result252[72]^and_result252[73]^and_result252[74]^and_result252[75]^and_result252[76]^and_result252[77]^and_result252[78]^and_result252[79]^and_result252[80]^and_result252[81]^and_result252[82]^and_result252[83]^and_result252[84]^and_result252[85]^and_result252[86]^and_result252[87]^and_result252[88]^and_result252[89]^and_result252[90]^and_result252[91]^and_result252[92]^and_result252[93]^and_result252[94]^and_result252[95]^and_result252[96]^and_result252[97]^and_result252[98]^and_result252[99]^and_result252[100]^and_result252[101]^and_result252[102]^and_result252[103]^and_result252[104]^and_result252[105]^and_result252[106]^and_result252[107]^and_result252[108]^and_result252[109]^and_result252[110]^and_result252[111]^and_result252[112]^and_result252[113]^and_result252[114]^and_result252[115]^and_result252[116]^and_result252[117]^and_result252[118]^and_result252[119]^and_result252[120]^and_result252[121]^and_result252[122]^and_result252[123]^and_result252[124]^and_result252[125]^and_result252[126]^and_result252[127]^and_result252[128]^and_result252[129]^and_result252[130]^and_result252[131]^and_result252[132]^and_result252[133]^and_result252[134]^and_result252[135]^and_result252[136]^and_result252[137]^and_result252[138]^and_result252[139]^and_result252[140]^and_result252[141]^and_result252[142]^and_result252[143]^and_result252[144]^and_result252[145]^and_result252[146]^and_result252[147]^and_result252[148]^and_result252[149]^and_result252[150]^and_result252[151]^and_result252[152]^and_result252[153]^and_result252[154]^and_result252[155]^and_result252[156]^and_result252[157]^and_result252[158]^and_result252[159]^and_result252[160]^and_result252[161]^and_result252[162]^and_result252[163]^and_result252[164]^and_result252[165]^and_result252[166]^and_result252[167]^and_result252[168]^and_result252[169]^and_result252[170]^and_result252[171]^and_result252[172]^and_result252[173]^and_result252[174]^and_result252[175]^and_result252[176]^and_result252[177]^and_result252[178]^and_result252[179]^and_result252[180]^and_result252[181]^and_result252[182]^and_result252[183]^and_result252[184]^and_result252[185]^and_result252[186]^and_result252[187]^and_result252[188]^and_result252[189]^and_result252[190]^and_result252[191]^and_result252[192]^and_result252[193]^and_result252[194]^and_result252[195]^and_result252[196]^and_result252[197]^and_result252[198]^and_result252[199]^and_result252[200]^and_result252[201]^and_result252[202]^and_result252[203]^and_result252[204]^and_result252[205]^and_result252[206]^and_result252[207]^and_result252[208]^and_result252[209]^and_result252[210]^and_result252[211]^and_result252[212]^and_result252[213]^and_result252[214]^and_result252[215]^and_result252[216]^and_result252[217]^and_result252[218]^and_result252[219]^and_result252[220]^and_result252[221]^and_result252[222]^and_result252[223]^and_result252[224]^and_result252[225]^and_result252[226]^and_result252[227]^and_result252[228]^and_result252[229]^and_result252[230]^and_result252[231]^and_result252[232]^and_result252[233]^and_result252[234]^and_result252[235]^and_result252[236]^and_result252[237]^and_result252[238]^and_result252[239]^and_result252[240]^and_result252[241]^and_result252[242]^and_result252[243]^and_result252[244]^and_result252[245]^and_result252[246]^and_result252[247]^and_result252[248]^and_result252[249]^and_result252[250]^and_result252[251]^and_result252[252]^and_result252[253]^and_result252[254];
assign key[253]=and_result253[0]^and_result253[1]^and_result253[2]^and_result253[3]^and_result253[4]^and_result253[5]^and_result253[6]^and_result253[7]^and_result253[8]^and_result253[9]^and_result253[10]^and_result253[11]^and_result253[12]^and_result253[13]^and_result253[14]^and_result253[15]^and_result253[16]^and_result253[17]^and_result253[18]^and_result253[19]^and_result253[20]^and_result253[21]^and_result253[22]^and_result253[23]^and_result253[24]^and_result253[25]^and_result253[26]^and_result253[27]^and_result253[28]^and_result253[29]^and_result253[30]^and_result253[31]^and_result253[32]^and_result253[33]^and_result253[34]^and_result253[35]^and_result253[36]^and_result253[37]^and_result253[38]^and_result253[39]^and_result253[40]^and_result253[41]^and_result253[42]^and_result253[43]^and_result253[44]^and_result253[45]^and_result253[46]^and_result253[47]^and_result253[48]^and_result253[49]^and_result253[50]^and_result253[51]^and_result253[52]^and_result253[53]^and_result253[54]^and_result253[55]^and_result253[56]^and_result253[57]^and_result253[58]^and_result253[59]^and_result253[60]^and_result253[61]^and_result253[62]^and_result253[63]^and_result253[64]^and_result253[65]^and_result253[66]^and_result253[67]^and_result253[68]^and_result253[69]^and_result253[70]^and_result253[71]^and_result253[72]^and_result253[73]^and_result253[74]^and_result253[75]^and_result253[76]^and_result253[77]^and_result253[78]^and_result253[79]^and_result253[80]^and_result253[81]^and_result253[82]^and_result253[83]^and_result253[84]^and_result253[85]^and_result253[86]^and_result253[87]^and_result253[88]^and_result253[89]^and_result253[90]^and_result253[91]^and_result253[92]^and_result253[93]^and_result253[94]^and_result253[95]^and_result253[96]^and_result253[97]^and_result253[98]^and_result253[99]^and_result253[100]^and_result253[101]^and_result253[102]^and_result253[103]^and_result253[104]^and_result253[105]^and_result253[106]^and_result253[107]^and_result253[108]^and_result253[109]^and_result253[110]^and_result253[111]^and_result253[112]^and_result253[113]^and_result253[114]^and_result253[115]^and_result253[116]^and_result253[117]^and_result253[118]^and_result253[119]^and_result253[120]^and_result253[121]^and_result253[122]^and_result253[123]^and_result253[124]^and_result253[125]^and_result253[126]^and_result253[127]^and_result253[128]^and_result253[129]^and_result253[130]^and_result253[131]^and_result253[132]^and_result253[133]^and_result253[134]^and_result253[135]^and_result253[136]^and_result253[137]^and_result253[138]^and_result253[139]^and_result253[140]^and_result253[141]^and_result253[142]^and_result253[143]^and_result253[144]^and_result253[145]^and_result253[146]^and_result253[147]^and_result253[148]^and_result253[149]^and_result253[150]^and_result253[151]^and_result253[152]^and_result253[153]^and_result253[154]^and_result253[155]^and_result253[156]^and_result253[157]^and_result253[158]^and_result253[159]^and_result253[160]^and_result253[161]^and_result253[162]^and_result253[163]^and_result253[164]^and_result253[165]^and_result253[166]^and_result253[167]^and_result253[168]^and_result253[169]^and_result253[170]^and_result253[171]^and_result253[172]^and_result253[173]^and_result253[174]^and_result253[175]^and_result253[176]^and_result253[177]^and_result253[178]^and_result253[179]^and_result253[180]^and_result253[181]^and_result253[182]^and_result253[183]^and_result253[184]^and_result253[185]^and_result253[186]^and_result253[187]^and_result253[188]^and_result253[189]^and_result253[190]^and_result253[191]^and_result253[192]^and_result253[193]^and_result253[194]^and_result253[195]^and_result253[196]^and_result253[197]^and_result253[198]^and_result253[199]^and_result253[200]^and_result253[201]^and_result253[202]^and_result253[203]^and_result253[204]^and_result253[205]^and_result253[206]^and_result253[207]^and_result253[208]^and_result253[209]^and_result253[210]^and_result253[211]^and_result253[212]^and_result253[213]^and_result253[214]^and_result253[215]^and_result253[216]^and_result253[217]^and_result253[218]^and_result253[219]^and_result253[220]^and_result253[221]^and_result253[222]^and_result253[223]^and_result253[224]^and_result253[225]^and_result253[226]^and_result253[227]^and_result253[228]^and_result253[229]^and_result253[230]^and_result253[231]^and_result253[232]^and_result253[233]^and_result253[234]^and_result253[235]^and_result253[236]^and_result253[237]^and_result253[238]^and_result253[239]^and_result253[240]^and_result253[241]^and_result253[242]^and_result253[243]^and_result253[244]^and_result253[245]^and_result253[246]^and_result253[247]^and_result253[248]^and_result253[249]^and_result253[250]^and_result253[251]^and_result253[252]^and_result253[253]^and_result253[254];
assign key[254]=and_result254[0]^and_result254[1]^and_result254[2]^and_result254[3]^and_result254[4]^and_result254[5]^and_result254[6]^and_result254[7]^and_result254[8]^and_result254[9]^and_result254[10]^and_result254[11]^and_result254[12]^and_result254[13]^and_result254[14]^and_result254[15]^and_result254[16]^and_result254[17]^and_result254[18]^and_result254[19]^and_result254[20]^and_result254[21]^and_result254[22]^and_result254[23]^and_result254[24]^and_result254[25]^and_result254[26]^and_result254[27]^and_result254[28]^and_result254[29]^and_result254[30]^and_result254[31]^and_result254[32]^and_result254[33]^and_result254[34]^and_result254[35]^and_result254[36]^and_result254[37]^and_result254[38]^and_result254[39]^and_result254[40]^and_result254[41]^and_result254[42]^and_result254[43]^and_result254[44]^and_result254[45]^and_result254[46]^and_result254[47]^and_result254[48]^and_result254[49]^and_result254[50]^and_result254[51]^and_result254[52]^and_result254[53]^and_result254[54]^and_result254[55]^and_result254[56]^and_result254[57]^and_result254[58]^and_result254[59]^and_result254[60]^and_result254[61]^and_result254[62]^and_result254[63]^and_result254[64]^and_result254[65]^and_result254[66]^and_result254[67]^and_result254[68]^and_result254[69]^and_result254[70]^and_result254[71]^and_result254[72]^and_result254[73]^and_result254[74]^and_result254[75]^and_result254[76]^and_result254[77]^and_result254[78]^and_result254[79]^and_result254[80]^and_result254[81]^and_result254[82]^and_result254[83]^and_result254[84]^and_result254[85]^and_result254[86]^and_result254[87]^and_result254[88]^and_result254[89]^and_result254[90]^and_result254[91]^and_result254[92]^and_result254[93]^and_result254[94]^and_result254[95]^and_result254[96]^and_result254[97]^and_result254[98]^and_result254[99]^and_result254[100]^and_result254[101]^and_result254[102]^and_result254[103]^and_result254[104]^and_result254[105]^and_result254[106]^and_result254[107]^and_result254[108]^and_result254[109]^and_result254[110]^and_result254[111]^and_result254[112]^and_result254[113]^and_result254[114]^and_result254[115]^and_result254[116]^and_result254[117]^and_result254[118]^and_result254[119]^and_result254[120]^and_result254[121]^and_result254[122]^and_result254[123]^and_result254[124]^and_result254[125]^and_result254[126]^and_result254[127]^and_result254[128]^and_result254[129]^and_result254[130]^and_result254[131]^and_result254[132]^and_result254[133]^and_result254[134]^and_result254[135]^and_result254[136]^and_result254[137]^and_result254[138]^and_result254[139]^and_result254[140]^and_result254[141]^and_result254[142]^and_result254[143]^and_result254[144]^and_result254[145]^and_result254[146]^and_result254[147]^and_result254[148]^and_result254[149]^and_result254[150]^and_result254[151]^and_result254[152]^and_result254[153]^and_result254[154]^and_result254[155]^and_result254[156]^and_result254[157]^and_result254[158]^and_result254[159]^and_result254[160]^and_result254[161]^and_result254[162]^and_result254[163]^and_result254[164]^and_result254[165]^and_result254[166]^and_result254[167]^and_result254[168]^and_result254[169]^and_result254[170]^and_result254[171]^and_result254[172]^and_result254[173]^and_result254[174]^and_result254[175]^and_result254[176]^and_result254[177]^and_result254[178]^and_result254[179]^and_result254[180]^and_result254[181]^and_result254[182]^and_result254[183]^and_result254[184]^and_result254[185]^and_result254[186]^and_result254[187]^and_result254[188]^and_result254[189]^and_result254[190]^and_result254[191]^and_result254[192]^and_result254[193]^and_result254[194]^and_result254[195]^and_result254[196]^and_result254[197]^and_result254[198]^and_result254[199]^and_result254[200]^and_result254[201]^and_result254[202]^and_result254[203]^and_result254[204]^and_result254[205]^and_result254[206]^and_result254[207]^and_result254[208]^and_result254[209]^and_result254[210]^and_result254[211]^and_result254[212]^and_result254[213]^and_result254[214]^and_result254[215]^and_result254[216]^and_result254[217]^and_result254[218]^and_result254[219]^and_result254[220]^and_result254[221]^and_result254[222]^and_result254[223]^and_result254[224]^and_result254[225]^and_result254[226]^and_result254[227]^and_result254[228]^and_result254[229]^and_result254[230]^and_result254[231]^and_result254[232]^and_result254[233]^and_result254[234]^and_result254[235]^and_result254[236]^and_result254[237]^and_result254[238]^and_result254[239]^and_result254[240]^and_result254[241]^and_result254[242]^and_result254[243]^and_result254[244]^and_result254[245]^and_result254[246]^and_result254[247]^and_result254[248]^and_result254[249]^and_result254[250]^and_result254[251]^and_result254[252]^and_result254[253]^and_result254[254];
    
endmodule

module tapes2tmp_shares(
    input [`tapesLength-1:0] tapes,
    input [10:0] pos,
    
    output [`state_mask_length-1:0] tmp_shares
);
    assign tmp_shares[15:0]={tapes[pos], tapes[pos+2295], tapes[pos+4590], tapes[pos+6885], tapes[pos+9180], tapes[pos+11475], tapes[pos+13770], tapes[pos+16065], tapes[pos+18360], tapes[pos+20655], tapes[pos+22950], tapes[pos+25245], tapes[pos+27540], tapes[pos+29835], tapes[pos+32130], tapes[pos+34425]};
    assign tmp_shares[31:16]={tapes[pos+1], tapes[pos+2296], tapes[pos+4591], tapes[pos+6886], tapes[pos+9181], tapes[pos+11476], tapes[pos+13771], tapes[pos+16066], tapes[pos+18361], tapes[pos+20656], tapes[pos+22951], tapes[pos+25246], tapes[pos+27541], tapes[pos+29836], tapes[pos+32131], tapes[pos+34426]};
    assign tmp_shares[47:32]={tapes[pos+2], tapes[pos+2297], tapes[pos+4592], tapes[pos+6887], tapes[pos+9182], tapes[pos+11477], tapes[pos+13772], tapes[pos+16067], tapes[pos+18362], tapes[pos+20657], tapes[pos+22952], tapes[pos+25247], tapes[pos+27542], tapes[pos+29837], tapes[pos+32132], tapes[pos+34427]};
    assign tmp_shares[63:48]={tapes[pos+3], tapes[pos+2298], tapes[pos+4593], tapes[pos+6888], tapes[pos+9183], tapes[pos+11478], tapes[pos+13773], tapes[pos+16068], tapes[pos+18363], tapes[pos+20658], tapes[pos+22953], tapes[pos+25248], tapes[pos+27543], tapes[pos+29838], tapes[pos+32133], tapes[pos+34428]};
    assign tmp_shares[79:64]={tapes[pos+4], tapes[pos+2299], tapes[pos+4594], tapes[pos+6889], tapes[pos+9184], tapes[pos+11479], tapes[pos+13774], tapes[pos+16069], tapes[pos+18364], tapes[pos+20659], tapes[pos+22954], tapes[pos+25249], tapes[pos+27544], tapes[pos+29839], tapes[pos+32134], tapes[pos+34429]};
    assign tmp_shares[95:80]={tapes[pos+5], tapes[pos+2300], tapes[pos+4595], tapes[pos+6890], tapes[pos+9185], tapes[pos+11480], tapes[pos+13775], tapes[pos+16070], tapes[pos+18365], tapes[pos+20660], tapes[pos+22955], tapes[pos+25250], tapes[pos+27545], tapes[pos+29840], tapes[pos+32135], tapes[pos+34430]};
    assign tmp_shares[111:96]={tapes[pos+6], tapes[pos+2301], tapes[pos+4596], tapes[pos+6891], tapes[pos+9186], tapes[pos+11481], tapes[pos+13776], tapes[pos+16071], tapes[pos+18366], tapes[pos+20661], tapes[pos+22956], tapes[pos+25251], tapes[pos+27546], tapes[pos+29841], tapes[pos+32136], tapes[pos+34431]};
    assign tmp_shares[127:112]={tapes[pos+7], tapes[pos+2302], tapes[pos+4597], tapes[pos+6892], tapes[pos+9187], tapes[pos+11482], tapes[pos+13777], tapes[pos+16072], tapes[pos+18367], tapes[pos+20662], tapes[pos+22957], tapes[pos+25252], tapes[pos+27547], tapes[pos+29842], tapes[pos+32137], tapes[pos+34432]};
    assign tmp_shares[143:128]={tapes[pos+8], tapes[pos+2303], tapes[pos+4598], tapes[pos+6893], tapes[pos+9188], tapes[pos+11483], tapes[pos+13778], tapes[pos+16073], tapes[pos+18368], tapes[pos+20663], tapes[pos+22958], tapes[pos+25253], tapes[pos+27548], tapes[pos+29843], tapes[pos+32138], tapes[pos+34433]};
    assign tmp_shares[159:144]={tapes[pos+9], tapes[pos+2304], tapes[pos+4599], tapes[pos+6894], tapes[pos+9189], tapes[pos+11484], tapes[pos+13779], tapes[pos+16074], tapes[pos+18369], tapes[pos+20664], tapes[pos+22959], tapes[pos+25254], tapes[pos+27549], tapes[pos+29844], tapes[pos+32139], tapes[pos+34434]};
    assign tmp_shares[175:160]={tapes[pos+10], tapes[pos+2305], tapes[pos+4600], tapes[pos+6895], tapes[pos+9190], tapes[pos+11485], tapes[pos+13780], tapes[pos+16075], tapes[pos+18370], tapes[pos+20665], tapes[pos+22960], tapes[pos+25255], tapes[pos+27550], tapes[pos+29845], tapes[pos+32140], tapes[pos+34435]};
    assign tmp_shares[191:176]={tapes[pos+11], tapes[pos+2306], tapes[pos+4601], tapes[pos+6896], tapes[pos+9191], tapes[pos+11486], tapes[pos+13781], tapes[pos+16076], tapes[pos+18371], tapes[pos+20666], tapes[pos+22961], tapes[pos+25256], tapes[pos+27551], tapes[pos+29846], tapes[pos+32141], tapes[pos+34436]};
    assign tmp_shares[207:192]={tapes[pos+12], tapes[pos+2307], tapes[pos+4602], tapes[pos+6897], tapes[pos+9192], tapes[pos+11487], tapes[pos+13782], tapes[pos+16077], tapes[pos+18372], tapes[pos+20667], tapes[pos+22962], tapes[pos+25257], tapes[pos+27552], tapes[pos+29847], tapes[pos+32142], tapes[pos+34437]};
    assign tmp_shares[223:208]={tapes[pos+13], tapes[pos+2308], tapes[pos+4603], tapes[pos+6898], tapes[pos+9193], tapes[pos+11488], tapes[pos+13783], tapes[pos+16078], tapes[pos+18373], tapes[pos+20668], tapes[pos+22963], tapes[pos+25258], tapes[pos+27553], tapes[pos+29848], tapes[pos+32143], tapes[pos+34438]};
    assign tmp_shares[239:224]={tapes[pos+14], tapes[pos+2309], tapes[pos+4604], tapes[pos+6899], tapes[pos+9194], tapes[pos+11489], tapes[pos+13784], tapes[pos+16079], tapes[pos+18374], tapes[pos+20669], tapes[pos+22964], tapes[pos+25259], tapes[pos+27554], tapes[pos+29849], tapes[pos+32144], tapes[pos+34439]};
    assign tmp_shares[255:240]={tapes[pos+15], tapes[pos+2310], tapes[pos+4605], tapes[pos+6900], tapes[pos+9195], tapes[pos+11490], tapes[pos+13785], tapes[pos+16080], tapes[pos+18375], tapes[pos+20670], tapes[pos+22965], tapes[pos+25260], tapes[pos+27555], tapes[pos+29850], tapes[pos+32145], tapes[pos+34440]};
    assign tmp_shares[271:256]={tapes[pos+16], tapes[pos+2311], tapes[pos+4606], tapes[pos+6901], tapes[pos+9196], tapes[pos+11491], tapes[pos+13786], tapes[pos+16081], tapes[pos+18376], tapes[pos+20671], tapes[pos+22966], tapes[pos+25261], tapes[pos+27556], tapes[pos+29851], tapes[pos+32146], tapes[pos+34441]};
    assign tmp_shares[287:272]={tapes[pos+17], tapes[pos+2312], tapes[pos+4607], tapes[pos+6902], tapes[pos+9197], tapes[pos+11492], tapes[pos+13787], tapes[pos+16082], tapes[pos+18377], tapes[pos+20672], tapes[pos+22967], tapes[pos+25262], tapes[pos+27557], tapes[pos+29852], tapes[pos+32147], tapes[pos+34442]};
    assign tmp_shares[303:288]={tapes[pos+18], tapes[pos+2313], tapes[pos+4608], tapes[pos+6903], tapes[pos+9198], tapes[pos+11493], tapes[pos+13788], tapes[pos+16083], tapes[pos+18378], tapes[pos+20673], tapes[pos+22968], tapes[pos+25263], tapes[pos+27558], tapes[pos+29853], tapes[pos+32148], tapes[pos+34443]};
    assign tmp_shares[319:304]={tapes[pos+19], tapes[pos+2314], tapes[pos+4609], tapes[pos+6904], tapes[pos+9199], tapes[pos+11494], tapes[pos+13789], tapes[pos+16084], tapes[pos+18379], tapes[pos+20674], tapes[pos+22969], tapes[pos+25264], tapes[pos+27559], tapes[pos+29854], tapes[pos+32149], tapes[pos+34444]};
    assign tmp_shares[335:320]={tapes[pos+20], tapes[pos+2315], tapes[pos+4610], tapes[pos+6905], tapes[pos+9200], tapes[pos+11495], tapes[pos+13790], tapes[pos+16085], tapes[pos+18380], tapes[pos+20675], tapes[pos+22970], tapes[pos+25265], tapes[pos+27560], tapes[pos+29855], tapes[pos+32150], tapes[pos+34445]};
    assign tmp_shares[351:336]={tapes[pos+21], tapes[pos+2316], tapes[pos+4611], tapes[pos+6906], tapes[pos+9201], tapes[pos+11496], tapes[pos+13791], tapes[pos+16086], tapes[pos+18381], tapes[pos+20676], tapes[pos+22971], tapes[pos+25266], tapes[pos+27561], tapes[pos+29856], tapes[pos+32151], tapes[pos+34446]};
    assign tmp_shares[367:352]={tapes[pos+22], tapes[pos+2317], tapes[pos+4612], tapes[pos+6907], tapes[pos+9202], tapes[pos+11497], tapes[pos+13792], tapes[pos+16087], tapes[pos+18382], tapes[pos+20677], tapes[pos+22972], tapes[pos+25267], tapes[pos+27562], tapes[pos+29857], tapes[pos+32152], tapes[pos+34447]};
    assign tmp_shares[383:368]={tapes[pos+23], tapes[pos+2318], tapes[pos+4613], tapes[pos+6908], tapes[pos+9203], tapes[pos+11498], tapes[pos+13793], tapes[pos+16088], tapes[pos+18383], tapes[pos+20678], tapes[pos+22973], tapes[pos+25268], tapes[pos+27563], tapes[pos+29858], tapes[pos+32153], tapes[pos+34448]};
    assign tmp_shares[399:384]={tapes[pos+24], tapes[pos+2319], tapes[pos+4614], tapes[pos+6909], tapes[pos+9204], tapes[pos+11499], tapes[pos+13794], tapes[pos+16089], tapes[pos+18384], tapes[pos+20679], tapes[pos+22974], tapes[pos+25269], tapes[pos+27564], tapes[pos+29859], tapes[pos+32154], tapes[pos+34449]};
    assign tmp_shares[415:400]={tapes[pos+25], tapes[pos+2320], tapes[pos+4615], tapes[pos+6910], tapes[pos+9205], tapes[pos+11500], tapes[pos+13795], tapes[pos+16090], tapes[pos+18385], tapes[pos+20680], tapes[pos+22975], tapes[pos+25270], tapes[pos+27565], tapes[pos+29860], tapes[pos+32155], tapes[pos+34450]};
    assign tmp_shares[431:416]={tapes[pos+26], tapes[pos+2321], tapes[pos+4616], tapes[pos+6911], tapes[pos+9206], tapes[pos+11501], tapes[pos+13796], tapes[pos+16091], tapes[pos+18386], tapes[pos+20681], tapes[pos+22976], tapes[pos+25271], tapes[pos+27566], tapes[pos+29861], tapes[pos+32156], tapes[pos+34451]};
    assign tmp_shares[447:432]={tapes[pos+27], tapes[pos+2322], tapes[pos+4617], tapes[pos+6912], tapes[pos+9207], tapes[pos+11502], tapes[pos+13797], tapes[pos+16092], tapes[pos+18387], tapes[pos+20682], tapes[pos+22977], tapes[pos+25272], tapes[pos+27567], tapes[pos+29862], tapes[pos+32157], tapes[pos+34452]};
    assign tmp_shares[463:448]={tapes[pos+28], tapes[pos+2323], tapes[pos+4618], tapes[pos+6913], tapes[pos+9208], tapes[pos+11503], tapes[pos+13798], tapes[pos+16093], tapes[pos+18388], tapes[pos+20683], tapes[pos+22978], tapes[pos+25273], tapes[pos+27568], tapes[pos+29863], tapes[pos+32158], tapes[pos+34453]};
    assign tmp_shares[479:464]={tapes[pos+29], tapes[pos+2324], tapes[pos+4619], tapes[pos+6914], tapes[pos+9209], tapes[pos+11504], tapes[pos+13799], tapes[pos+16094], tapes[pos+18389], tapes[pos+20684], tapes[pos+22979], tapes[pos+25274], tapes[pos+27569], tapes[pos+29864], tapes[pos+32159], tapes[pos+34454]};
    assign tmp_shares[495:480]={tapes[pos+30], tapes[pos+2325], tapes[pos+4620], tapes[pos+6915], tapes[pos+9210], tapes[pos+11505], tapes[pos+13800], tapes[pos+16095], tapes[pos+18390], tapes[pos+20685], tapes[pos+22980], tapes[pos+25275], tapes[pos+27570], tapes[pos+29865], tapes[pos+32160], tapes[pos+34455]};
    assign tmp_shares[511:496]={tapes[pos+31], tapes[pos+2326], tapes[pos+4621], tapes[pos+6916], tapes[pos+9211], tapes[pos+11506], tapes[pos+13801], tapes[pos+16096], tapes[pos+18391], tapes[pos+20686], tapes[pos+22981], tapes[pos+25276], tapes[pos+27571], tapes[pos+29866], tapes[pos+32161], tapes[pos+34456]};
    assign tmp_shares[527:512]={tapes[pos+32], tapes[pos+2327], tapes[pos+4622], tapes[pos+6917], tapes[pos+9212], tapes[pos+11507], tapes[pos+13802], tapes[pos+16097], tapes[pos+18392], tapes[pos+20687], tapes[pos+22982], tapes[pos+25277], tapes[pos+27572], tapes[pos+29867], tapes[pos+32162], tapes[pos+34457]};
    assign tmp_shares[543:528]={tapes[pos+33], tapes[pos+2328], tapes[pos+4623], tapes[pos+6918], tapes[pos+9213], tapes[pos+11508], tapes[pos+13803], tapes[pos+16098], tapes[pos+18393], tapes[pos+20688], tapes[pos+22983], tapes[pos+25278], tapes[pos+27573], tapes[pos+29868], tapes[pos+32163], tapes[pos+34458]};
    assign tmp_shares[559:544]={tapes[pos+34], tapes[pos+2329], tapes[pos+4624], tapes[pos+6919], tapes[pos+9214], tapes[pos+11509], tapes[pos+13804], tapes[pos+16099], tapes[pos+18394], tapes[pos+20689], tapes[pos+22984], tapes[pos+25279], tapes[pos+27574], tapes[pos+29869], tapes[pos+32164], tapes[pos+34459]};
    assign tmp_shares[575:560]={tapes[pos+35], tapes[pos+2330], tapes[pos+4625], tapes[pos+6920], tapes[pos+9215], tapes[pos+11510], tapes[pos+13805], tapes[pos+16100], tapes[pos+18395], tapes[pos+20690], tapes[pos+22985], tapes[pos+25280], tapes[pos+27575], tapes[pos+29870], tapes[pos+32165], tapes[pos+34460]};
    assign tmp_shares[591:576]={tapes[pos+36], tapes[pos+2331], tapes[pos+4626], tapes[pos+6921], tapes[pos+9216], tapes[pos+11511], tapes[pos+13806], tapes[pos+16101], tapes[pos+18396], tapes[pos+20691], tapes[pos+22986], tapes[pos+25281], tapes[pos+27576], tapes[pos+29871], tapes[pos+32166], tapes[pos+34461]};
    assign tmp_shares[607:592]={tapes[pos+37], tapes[pos+2332], tapes[pos+4627], tapes[pos+6922], tapes[pos+9217], tapes[pos+11512], tapes[pos+13807], tapes[pos+16102], tapes[pos+18397], tapes[pos+20692], tapes[pos+22987], tapes[pos+25282], tapes[pos+27577], tapes[pos+29872], tapes[pos+32167], tapes[pos+34462]};
    assign tmp_shares[623:608]={tapes[pos+38], tapes[pos+2333], tapes[pos+4628], tapes[pos+6923], tapes[pos+9218], tapes[pos+11513], tapes[pos+13808], tapes[pos+16103], tapes[pos+18398], tapes[pos+20693], tapes[pos+22988], tapes[pos+25283], tapes[pos+27578], tapes[pos+29873], tapes[pos+32168], tapes[pos+34463]};
    assign tmp_shares[639:624]={tapes[pos+39], tapes[pos+2334], tapes[pos+4629], tapes[pos+6924], tapes[pos+9219], tapes[pos+11514], tapes[pos+13809], tapes[pos+16104], tapes[pos+18399], tapes[pos+20694], tapes[pos+22989], tapes[pos+25284], tapes[pos+27579], tapes[pos+29874], tapes[pos+32169], tapes[pos+34464]};
    assign tmp_shares[655:640]={tapes[pos+40], tapes[pos+2335], tapes[pos+4630], tapes[pos+6925], tapes[pos+9220], tapes[pos+11515], tapes[pos+13810], tapes[pos+16105], tapes[pos+18400], tapes[pos+20695], tapes[pos+22990], tapes[pos+25285], tapes[pos+27580], tapes[pos+29875], tapes[pos+32170], tapes[pos+34465]};
    assign tmp_shares[671:656]={tapes[pos+41], tapes[pos+2336], tapes[pos+4631], tapes[pos+6926], tapes[pos+9221], tapes[pos+11516], tapes[pos+13811], tapes[pos+16106], tapes[pos+18401], tapes[pos+20696], tapes[pos+22991], tapes[pos+25286], tapes[pos+27581], tapes[pos+29876], tapes[pos+32171], tapes[pos+34466]};
    assign tmp_shares[687:672]={tapes[pos+42], tapes[pos+2337], tapes[pos+4632], tapes[pos+6927], tapes[pos+9222], tapes[pos+11517], tapes[pos+13812], tapes[pos+16107], tapes[pos+18402], tapes[pos+20697], tapes[pos+22992], tapes[pos+25287], tapes[pos+27582], tapes[pos+29877], tapes[pos+32172], tapes[pos+34467]};
    assign tmp_shares[703:688]={tapes[pos+43], tapes[pos+2338], tapes[pos+4633], tapes[pos+6928], tapes[pos+9223], tapes[pos+11518], tapes[pos+13813], tapes[pos+16108], tapes[pos+18403], tapes[pos+20698], tapes[pos+22993], tapes[pos+25288], tapes[pos+27583], tapes[pos+29878], tapes[pos+32173], tapes[pos+34468]};
    assign tmp_shares[719:704]={tapes[pos+44], tapes[pos+2339], tapes[pos+4634], tapes[pos+6929], tapes[pos+9224], tapes[pos+11519], tapes[pos+13814], tapes[pos+16109], tapes[pos+18404], tapes[pos+20699], tapes[pos+22994], tapes[pos+25289], tapes[pos+27584], tapes[pos+29879], tapes[pos+32174], tapes[pos+34469]};
    assign tmp_shares[735:720]={tapes[pos+45], tapes[pos+2340], tapes[pos+4635], tapes[pos+6930], tapes[pos+9225], tapes[pos+11520], tapes[pos+13815], tapes[pos+16110], tapes[pos+18405], tapes[pos+20700], tapes[pos+22995], tapes[pos+25290], tapes[pos+27585], tapes[pos+29880], tapes[pos+32175], tapes[pos+34470]};
    assign tmp_shares[751:736]={tapes[pos+46], tapes[pos+2341], tapes[pos+4636], tapes[pos+6931], tapes[pos+9226], tapes[pos+11521], tapes[pos+13816], tapes[pos+16111], tapes[pos+18406], tapes[pos+20701], tapes[pos+22996], tapes[pos+25291], tapes[pos+27586], tapes[pos+29881], tapes[pos+32176], tapes[pos+34471]};
    assign tmp_shares[767:752]={tapes[pos+47], tapes[pos+2342], tapes[pos+4637], tapes[pos+6932], tapes[pos+9227], tapes[pos+11522], tapes[pos+13817], tapes[pos+16112], tapes[pos+18407], tapes[pos+20702], tapes[pos+22997], tapes[pos+25292], tapes[pos+27587], tapes[pos+29882], tapes[pos+32177], tapes[pos+34472]};
    assign tmp_shares[783:768]={tapes[pos+48], tapes[pos+2343], tapes[pos+4638], tapes[pos+6933], tapes[pos+9228], tapes[pos+11523], tapes[pos+13818], tapes[pos+16113], tapes[pos+18408], tapes[pos+20703], tapes[pos+22998], tapes[pos+25293], tapes[pos+27588], tapes[pos+29883], tapes[pos+32178], tapes[pos+34473]};
    assign tmp_shares[799:784]={tapes[pos+49], tapes[pos+2344], tapes[pos+4639], tapes[pos+6934], tapes[pos+9229], tapes[pos+11524], tapes[pos+13819], tapes[pos+16114], tapes[pos+18409], tapes[pos+20704], tapes[pos+22999], tapes[pos+25294], tapes[pos+27589], tapes[pos+29884], tapes[pos+32179], tapes[pos+34474]};
    assign tmp_shares[815:800]={tapes[pos+50], tapes[pos+2345], tapes[pos+4640], tapes[pos+6935], tapes[pos+9230], tapes[pos+11525], tapes[pos+13820], tapes[pos+16115], tapes[pos+18410], tapes[pos+20705], tapes[pos+23000], tapes[pos+25295], tapes[pos+27590], tapes[pos+29885], tapes[pos+32180], tapes[pos+34475]};
    assign tmp_shares[831:816]={tapes[pos+51], tapes[pos+2346], tapes[pos+4641], tapes[pos+6936], tapes[pos+9231], tapes[pos+11526], tapes[pos+13821], tapes[pos+16116], tapes[pos+18411], tapes[pos+20706], tapes[pos+23001], tapes[pos+25296], tapes[pos+27591], tapes[pos+29886], tapes[pos+32181], tapes[pos+34476]};
    assign tmp_shares[847:832]={tapes[pos+52], tapes[pos+2347], tapes[pos+4642], tapes[pos+6937], tapes[pos+9232], tapes[pos+11527], tapes[pos+13822], tapes[pos+16117], tapes[pos+18412], tapes[pos+20707], tapes[pos+23002], tapes[pos+25297], tapes[pos+27592], tapes[pos+29887], tapes[pos+32182], tapes[pos+34477]};
    assign tmp_shares[863:848]={tapes[pos+53], tapes[pos+2348], tapes[pos+4643], tapes[pos+6938], tapes[pos+9233], tapes[pos+11528], tapes[pos+13823], tapes[pos+16118], tapes[pos+18413], tapes[pos+20708], tapes[pos+23003], tapes[pos+25298], tapes[pos+27593], tapes[pos+29888], tapes[pos+32183], tapes[pos+34478]};
    assign tmp_shares[879:864]={tapes[pos+54], tapes[pos+2349], tapes[pos+4644], tapes[pos+6939], tapes[pos+9234], tapes[pos+11529], tapes[pos+13824], tapes[pos+16119], tapes[pos+18414], tapes[pos+20709], tapes[pos+23004], tapes[pos+25299], tapes[pos+27594], tapes[pos+29889], tapes[pos+32184], tapes[pos+34479]};
    assign tmp_shares[895:880]={tapes[pos+55], tapes[pos+2350], tapes[pos+4645], tapes[pos+6940], tapes[pos+9235], tapes[pos+11530], tapes[pos+13825], tapes[pos+16120], tapes[pos+18415], tapes[pos+20710], tapes[pos+23005], tapes[pos+25300], tapes[pos+27595], tapes[pos+29890], tapes[pos+32185], tapes[pos+34480]};
    assign tmp_shares[911:896]={tapes[pos+56], tapes[pos+2351], tapes[pos+4646], tapes[pos+6941], tapes[pos+9236], tapes[pos+11531], tapes[pos+13826], tapes[pos+16121], tapes[pos+18416], tapes[pos+20711], tapes[pos+23006], tapes[pos+25301], tapes[pos+27596], tapes[pos+29891], tapes[pos+32186], tapes[pos+34481]};
    assign tmp_shares[927:912]={tapes[pos+57], tapes[pos+2352], tapes[pos+4647], tapes[pos+6942], tapes[pos+9237], tapes[pos+11532], tapes[pos+13827], tapes[pos+16122], tapes[pos+18417], tapes[pos+20712], tapes[pos+23007], tapes[pos+25302], tapes[pos+27597], tapes[pos+29892], tapes[pos+32187], tapes[pos+34482]};
    assign tmp_shares[943:928]={tapes[pos+58], tapes[pos+2353], tapes[pos+4648], tapes[pos+6943], tapes[pos+9238], tapes[pos+11533], tapes[pos+13828], tapes[pos+16123], tapes[pos+18418], tapes[pos+20713], tapes[pos+23008], tapes[pos+25303], tapes[pos+27598], tapes[pos+29893], tapes[pos+32188], tapes[pos+34483]};
    assign tmp_shares[959:944]={tapes[pos+59], tapes[pos+2354], tapes[pos+4649], tapes[pos+6944], tapes[pos+9239], tapes[pos+11534], tapes[pos+13829], tapes[pos+16124], tapes[pos+18419], tapes[pos+20714], tapes[pos+23009], tapes[pos+25304], tapes[pos+27599], tapes[pos+29894], tapes[pos+32189], tapes[pos+34484]};
    assign tmp_shares[975:960]={tapes[pos+60], tapes[pos+2355], tapes[pos+4650], tapes[pos+6945], tapes[pos+9240], tapes[pos+11535], tapes[pos+13830], tapes[pos+16125], tapes[pos+18420], tapes[pos+20715], tapes[pos+23010], tapes[pos+25305], tapes[pos+27600], tapes[pos+29895], tapes[pos+32190], tapes[pos+34485]};
    assign tmp_shares[991:976]={tapes[pos+61], tapes[pos+2356], tapes[pos+4651], tapes[pos+6946], tapes[pos+9241], tapes[pos+11536], tapes[pos+13831], tapes[pos+16126], tapes[pos+18421], tapes[pos+20716], tapes[pos+23011], tapes[pos+25306], tapes[pos+27601], tapes[pos+29896], tapes[pos+32191], tapes[pos+34486]};
    assign tmp_shares[1007:992]={tapes[pos+62], tapes[pos+2357], tapes[pos+4652], tapes[pos+6947], tapes[pos+9242], tapes[pos+11537], tapes[pos+13832], tapes[pos+16127], tapes[pos+18422], tapes[pos+20717], tapes[pos+23012], tapes[pos+25307], tapes[pos+27602], tapes[pos+29897], tapes[pos+32192], tapes[pos+34487]};
    assign tmp_shares[1023:1008]={tapes[pos+63], tapes[pos+2358], tapes[pos+4653], tapes[pos+6948], tapes[pos+9243], tapes[pos+11538], tapes[pos+13833], tapes[pos+16128], tapes[pos+18423], tapes[pos+20718], tapes[pos+23013], tapes[pos+25308], tapes[pos+27603], tapes[pos+29898], tapes[pos+32193], tapes[pos+34488]};
    assign tmp_shares[1039:1024]={tapes[pos+64], tapes[pos+2359], tapes[pos+4654], tapes[pos+6949], tapes[pos+9244], tapes[pos+11539], tapes[pos+13834], tapes[pos+16129], tapes[pos+18424], tapes[pos+20719], tapes[pos+23014], tapes[pos+25309], tapes[pos+27604], tapes[pos+29899], tapes[pos+32194], tapes[pos+34489]};
    assign tmp_shares[1055:1040]={tapes[pos+65], tapes[pos+2360], tapes[pos+4655], tapes[pos+6950], tapes[pos+9245], tapes[pos+11540], tapes[pos+13835], tapes[pos+16130], tapes[pos+18425], tapes[pos+20720], tapes[pos+23015], tapes[pos+25310], tapes[pos+27605], tapes[pos+29900], tapes[pos+32195], tapes[pos+34490]};
    assign tmp_shares[1071:1056]={tapes[pos+66], tapes[pos+2361], tapes[pos+4656], tapes[pos+6951], tapes[pos+9246], tapes[pos+11541], tapes[pos+13836], tapes[pos+16131], tapes[pos+18426], tapes[pos+20721], tapes[pos+23016], tapes[pos+25311], tapes[pos+27606], tapes[pos+29901], tapes[pos+32196], tapes[pos+34491]};
    assign tmp_shares[1087:1072]={tapes[pos+67], tapes[pos+2362], tapes[pos+4657], tapes[pos+6952], tapes[pos+9247], tapes[pos+11542], tapes[pos+13837], tapes[pos+16132], tapes[pos+18427], tapes[pos+20722], tapes[pos+23017], tapes[pos+25312], tapes[pos+27607], tapes[pos+29902], tapes[pos+32197], tapes[pos+34492]};
    assign tmp_shares[1103:1088]={tapes[pos+68], tapes[pos+2363], tapes[pos+4658], tapes[pos+6953], tapes[pos+9248], tapes[pos+11543], tapes[pos+13838], tapes[pos+16133], tapes[pos+18428], tapes[pos+20723], tapes[pos+23018], tapes[pos+25313], tapes[pos+27608], tapes[pos+29903], tapes[pos+32198], tapes[pos+34493]};
    assign tmp_shares[1119:1104]={tapes[pos+69], tapes[pos+2364], tapes[pos+4659], tapes[pos+6954], tapes[pos+9249], tapes[pos+11544], tapes[pos+13839], tapes[pos+16134], tapes[pos+18429], tapes[pos+20724], tapes[pos+23019], tapes[pos+25314], tapes[pos+27609], tapes[pos+29904], tapes[pos+32199], tapes[pos+34494]};
    assign tmp_shares[1135:1120]={tapes[pos+70], tapes[pos+2365], tapes[pos+4660], tapes[pos+6955], tapes[pos+9250], tapes[pos+11545], tapes[pos+13840], tapes[pos+16135], tapes[pos+18430], tapes[pos+20725], tapes[pos+23020], tapes[pos+25315], tapes[pos+27610], tapes[pos+29905], tapes[pos+32200], tapes[pos+34495]};
    assign tmp_shares[1151:1136]={tapes[pos+71], tapes[pos+2366], tapes[pos+4661], tapes[pos+6956], tapes[pos+9251], tapes[pos+11546], tapes[pos+13841], tapes[pos+16136], tapes[pos+18431], tapes[pos+20726], tapes[pos+23021], tapes[pos+25316], tapes[pos+27611], tapes[pos+29906], tapes[pos+32201], tapes[pos+34496]};
    assign tmp_shares[1167:1152]={tapes[pos+72], tapes[pos+2367], tapes[pos+4662], tapes[pos+6957], tapes[pos+9252], tapes[pos+11547], tapes[pos+13842], tapes[pos+16137], tapes[pos+18432], tapes[pos+20727], tapes[pos+23022], tapes[pos+25317], tapes[pos+27612], tapes[pos+29907], tapes[pos+32202], tapes[pos+34497]};
    assign tmp_shares[1183:1168]={tapes[pos+73], tapes[pos+2368], tapes[pos+4663], tapes[pos+6958], tapes[pos+9253], tapes[pos+11548], tapes[pos+13843], tapes[pos+16138], tapes[pos+18433], tapes[pos+20728], tapes[pos+23023], tapes[pos+25318], tapes[pos+27613], tapes[pos+29908], tapes[pos+32203], tapes[pos+34498]};
    assign tmp_shares[1199:1184]={tapes[pos+74], tapes[pos+2369], tapes[pos+4664], tapes[pos+6959], tapes[pos+9254], tapes[pos+11549], tapes[pos+13844], tapes[pos+16139], tapes[pos+18434], tapes[pos+20729], tapes[pos+23024], tapes[pos+25319], tapes[pos+27614], tapes[pos+29909], tapes[pos+32204], tapes[pos+34499]};
    assign tmp_shares[1215:1200]={tapes[pos+75], tapes[pos+2370], tapes[pos+4665], tapes[pos+6960], tapes[pos+9255], tapes[pos+11550], tapes[pos+13845], tapes[pos+16140], tapes[pos+18435], tapes[pos+20730], tapes[pos+23025], tapes[pos+25320], tapes[pos+27615], tapes[pos+29910], tapes[pos+32205], tapes[pos+34500]};
    assign tmp_shares[1231:1216]={tapes[pos+76], tapes[pos+2371], tapes[pos+4666], tapes[pos+6961], tapes[pos+9256], tapes[pos+11551], tapes[pos+13846], tapes[pos+16141], tapes[pos+18436], tapes[pos+20731], tapes[pos+23026], tapes[pos+25321], tapes[pos+27616], tapes[pos+29911], tapes[pos+32206], tapes[pos+34501]};
    assign tmp_shares[1247:1232]={tapes[pos+77], tapes[pos+2372], tapes[pos+4667], tapes[pos+6962], tapes[pos+9257], tapes[pos+11552], tapes[pos+13847], tapes[pos+16142], tapes[pos+18437], tapes[pos+20732], tapes[pos+23027], tapes[pos+25322], tapes[pos+27617], tapes[pos+29912], tapes[pos+32207], tapes[pos+34502]};
    assign tmp_shares[1263:1248]={tapes[pos+78], tapes[pos+2373], tapes[pos+4668], tapes[pos+6963], tapes[pos+9258], tapes[pos+11553], tapes[pos+13848], tapes[pos+16143], tapes[pos+18438], tapes[pos+20733], tapes[pos+23028], tapes[pos+25323], tapes[pos+27618], tapes[pos+29913], tapes[pos+32208], tapes[pos+34503]};
    assign tmp_shares[1279:1264]={tapes[pos+79], tapes[pos+2374], tapes[pos+4669], tapes[pos+6964], tapes[pos+9259], tapes[pos+11554], tapes[pos+13849], tapes[pos+16144], tapes[pos+18439], tapes[pos+20734], tapes[pos+23029], tapes[pos+25324], tapes[pos+27619], tapes[pos+29914], tapes[pos+32209], tapes[pos+34504]};
    assign tmp_shares[1295:1280]={tapes[pos+80], tapes[pos+2375], tapes[pos+4670], tapes[pos+6965], tapes[pos+9260], tapes[pos+11555], tapes[pos+13850], tapes[pos+16145], tapes[pos+18440], tapes[pos+20735], tapes[pos+23030], tapes[pos+25325], tapes[pos+27620], tapes[pos+29915], tapes[pos+32210], tapes[pos+34505]};
    assign tmp_shares[1311:1296]={tapes[pos+81], tapes[pos+2376], tapes[pos+4671], tapes[pos+6966], tapes[pos+9261], tapes[pos+11556], tapes[pos+13851], tapes[pos+16146], tapes[pos+18441], tapes[pos+20736], tapes[pos+23031], tapes[pos+25326], tapes[pos+27621], tapes[pos+29916], tapes[pos+32211], tapes[pos+34506]};
    assign tmp_shares[1327:1312]={tapes[pos+82], tapes[pos+2377], tapes[pos+4672], tapes[pos+6967], tapes[pos+9262], tapes[pos+11557], tapes[pos+13852], tapes[pos+16147], tapes[pos+18442], tapes[pos+20737], tapes[pos+23032], tapes[pos+25327], tapes[pos+27622], tapes[pos+29917], tapes[pos+32212], tapes[pos+34507]};
    assign tmp_shares[1343:1328]={tapes[pos+83], tapes[pos+2378], tapes[pos+4673], tapes[pos+6968], tapes[pos+9263], tapes[pos+11558], tapes[pos+13853], tapes[pos+16148], tapes[pos+18443], tapes[pos+20738], tapes[pos+23033], tapes[pos+25328], tapes[pos+27623], tapes[pos+29918], tapes[pos+32213], tapes[pos+34508]};
    assign tmp_shares[1359:1344]={tapes[pos+84], tapes[pos+2379], tapes[pos+4674], tapes[pos+6969], tapes[pos+9264], tapes[pos+11559], tapes[pos+13854], tapes[pos+16149], tapes[pos+18444], tapes[pos+20739], tapes[pos+23034], tapes[pos+25329], tapes[pos+27624], tapes[pos+29919], tapes[pos+32214], tapes[pos+34509]};
    assign tmp_shares[1375:1360]={tapes[pos+85], tapes[pos+2380], tapes[pos+4675], tapes[pos+6970], tapes[pos+9265], tapes[pos+11560], tapes[pos+13855], tapes[pos+16150], tapes[pos+18445], tapes[pos+20740], tapes[pos+23035], tapes[pos+25330], tapes[pos+27625], tapes[pos+29920], tapes[pos+32215], tapes[pos+34510]};
    assign tmp_shares[1391:1376]={tapes[pos+86], tapes[pos+2381], tapes[pos+4676], tapes[pos+6971], tapes[pos+9266], tapes[pos+11561], tapes[pos+13856], tapes[pos+16151], tapes[pos+18446], tapes[pos+20741], tapes[pos+23036], tapes[pos+25331], tapes[pos+27626], tapes[pos+29921], tapes[pos+32216], tapes[pos+34511]};
    assign tmp_shares[1407:1392]={tapes[pos+87], tapes[pos+2382], tapes[pos+4677], tapes[pos+6972], tapes[pos+9267], tapes[pos+11562], tapes[pos+13857], tapes[pos+16152], tapes[pos+18447], tapes[pos+20742], tapes[pos+23037], tapes[pos+25332], tapes[pos+27627], tapes[pos+29922], tapes[pos+32217], tapes[pos+34512]};
    assign tmp_shares[1423:1408]={tapes[pos+88], tapes[pos+2383], tapes[pos+4678], tapes[pos+6973], tapes[pos+9268], tapes[pos+11563], tapes[pos+13858], tapes[pos+16153], tapes[pos+18448], tapes[pos+20743], tapes[pos+23038], tapes[pos+25333], tapes[pos+27628], tapes[pos+29923], tapes[pos+32218], tapes[pos+34513]};
    assign tmp_shares[1439:1424]={tapes[pos+89], tapes[pos+2384], tapes[pos+4679], tapes[pos+6974], tapes[pos+9269], tapes[pos+11564], tapes[pos+13859], tapes[pos+16154], tapes[pos+18449], tapes[pos+20744], tapes[pos+23039], tapes[pos+25334], tapes[pos+27629], tapes[pos+29924], tapes[pos+32219], tapes[pos+34514]};
    assign tmp_shares[1455:1440]={tapes[pos+90], tapes[pos+2385], tapes[pos+4680], tapes[pos+6975], tapes[pos+9270], tapes[pos+11565], tapes[pos+13860], tapes[pos+16155], tapes[pos+18450], tapes[pos+20745], tapes[pos+23040], tapes[pos+25335], tapes[pos+27630], tapes[pos+29925], tapes[pos+32220], tapes[pos+34515]};
    assign tmp_shares[1471:1456]={tapes[pos+91], tapes[pos+2386], tapes[pos+4681], tapes[pos+6976], tapes[pos+9271], tapes[pos+11566], tapes[pos+13861], tapes[pos+16156], tapes[pos+18451], tapes[pos+20746], tapes[pos+23041], tapes[pos+25336], tapes[pos+27631], tapes[pos+29926], tapes[pos+32221], tapes[pos+34516]};
    assign tmp_shares[1487:1472]={tapes[pos+92], tapes[pos+2387], tapes[pos+4682], tapes[pos+6977], tapes[pos+9272], tapes[pos+11567], tapes[pos+13862], tapes[pos+16157], tapes[pos+18452], tapes[pos+20747], tapes[pos+23042], tapes[pos+25337], tapes[pos+27632], tapes[pos+29927], tapes[pos+32222], tapes[pos+34517]};
    assign tmp_shares[1503:1488]={tapes[pos+93], tapes[pos+2388], tapes[pos+4683], tapes[pos+6978], tapes[pos+9273], tapes[pos+11568], tapes[pos+13863], tapes[pos+16158], tapes[pos+18453], tapes[pos+20748], tapes[pos+23043], tapes[pos+25338], tapes[pos+27633], tapes[pos+29928], tapes[pos+32223], tapes[pos+34518]};
    assign tmp_shares[1519:1504]={tapes[pos+94], tapes[pos+2389], tapes[pos+4684], tapes[pos+6979], tapes[pos+9274], tapes[pos+11569], tapes[pos+13864], tapes[pos+16159], tapes[pos+18454], tapes[pos+20749], tapes[pos+23044], tapes[pos+25339], tapes[pos+27634], tapes[pos+29929], tapes[pos+32224], tapes[pos+34519]};
    assign tmp_shares[1535:1520]={tapes[pos+95], tapes[pos+2390], tapes[pos+4685], tapes[pos+6980], tapes[pos+9275], tapes[pos+11570], tapes[pos+13865], tapes[pos+16160], tapes[pos+18455], tapes[pos+20750], tapes[pos+23045], tapes[pos+25340], tapes[pos+27635], tapes[pos+29930], tapes[pos+32225], tapes[pos+34520]};
    assign tmp_shares[1551:1536]={tapes[pos+96], tapes[pos+2391], tapes[pos+4686], tapes[pos+6981], tapes[pos+9276], tapes[pos+11571], tapes[pos+13866], tapes[pos+16161], tapes[pos+18456], tapes[pos+20751], tapes[pos+23046], tapes[pos+25341], tapes[pos+27636], tapes[pos+29931], tapes[pos+32226], tapes[pos+34521]};
    assign tmp_shares[1567:1552]={tapes[pos+97], tapes[pos+2392], tapes[pos+4687], tapes[pos+6982], tapes[pos+9277], tapes[pos+11572], tapes[pos+13867], tapes[pos+16162], tapes[pos+18457], tapes[pos+20752], tapes[pos+23047], tapes[pos+25342], tapes[pos+27637], tapes[pos+29932], tapes[pos+32227], tapes[pos+34522]};
    assign tmp_shares[1583:1568]={tapes[pos+98], tapes[pos+2393], tapes[pos+4688], tapes[pos+6983], tapes[pos+9278], tapes[pos+11573], tapes[pos+13868], tapes[pos+16163], tapes[pos+18458], tapes[pos+20753], tapes[pos+23048], tapes[pos+25343], tapes[pos+27638], tapes[pos+29933], tapes[pos+32228], tapes[pos+34523]};
    assign tmp_shares[1599:1584]={tapes[pos+99], tapes[pos+2394], tapes[pos+4689], tapes[pos+6984], tapes[pos+9279], tapes[pos+11574], tapes[pos+13869], tapes[pos+16164], tapes[pos+18459], tapes[pos+20754], tapes[pos+23049], tapes[pos+25344], tapes[pos+27639], tapes[pos+29934], tapes[pos+32229], tapes[pos+34524]};
    assign tmp_shares[1615:1600]={tapes[pos+100], tapes[pos+2395], tapes[pos+4690], tapes[pos+6985], tapes[pos+9280], tapes[pos+11575], tapes[pos+13870], tapes[pos+16165], tapes[pos+18460], tapes[pos+20755], tapes[pos+23050], tapes[pos+25345], tapes[pos+27640], tapes[pos+29935], tapes[pos+32230], tapes[pos+34525]};
    assign tmp_shares[1631:1616]={tapes[pos+101], tapes[pos+2396], tapes[pos+4691], tapes[pos+6986], tapes[pos+9281], tapes[pos+11576], tapes[pos+13871], tapes[pos+16166], tapes[pos+18461], tapes[pos+20756], tapes[pos+23051], tapes[pos+25346], tapes[pos+27641], tapes[pos+29936], tapes[pos+32231], tapes[pos+34526]};
    assign tmp_shares[1647:1632]={tapes[pos+102], tapes[pos+2397], tapes[pos+4692], tapes[pos+6987], tapes[pos+9282], tapes[pos+11577], tapes[pos+13872], tapes[pos+16167], tapes[pos+18462], tapes[pos+20757], tapes[pos+23052], tapes[pos+25347], tapes[pos+27642], tapes[pos+29937], tapes[pos+32232], tapes[pos+34527]};
    assign tmp_shares[1663:1648]={tapes[pos+103], tapes[pos+2398], tapes[pos+4693], tapes[pos+6988], tapes[pos+9283], tapes[pos+11578], tapes[pos+13873], tapes[pos+16168], tapes[pos+18463], tapes[pos+20758], tapes[pos+23053], tapes[pos+25348], tapes[pos+27643], tapes[pos+29938], tapes[pos+32233], tapes[pos+34528]};
    assign tmp_shares[1679:1664]={tapes[pos+104], tapes[pos+2399], tapes[pos+4694], tapes[pos+6989], tapes[pos+9284], tapes[pos+11579], tapes[pos+13874], tapes[pos+16169], tapes[pos+18464], tapes[pos+20759], tapes[pos+23054], tapes[pos+25349], tapes[pos+27644], tapes[pos+29939], tapes[pos+32234], tapes[pos+34529]};
    assign tmp_shares[1695:1680]={tapes[pos+105], tapes[pos+2400], tapes[pos+4695], tapes[pos+6990], tapes[pos+9285], tapes[pos+11580], tapes[pos+13875], tapes[pos+16170], tapes[pos+18465], tapes[pos+20760], tapes[pos+23055], tapes[pos+25350], tapes[pos+27645], tapes[pos+29940], tapes[pos+32235], tapes[pos+34530]};
    assign tmp_shares[1711:1696]={tapes[pos+106], tapes[pos+2401], tapes[pos+4696], tapes[pos+6991], tapes[pos+9286], tapes[pos+11581], tapes[pos+13876], tapes[pos+16171], tapes[pos+18466], tapes[pos+20761], tapes[pos+23056], tapes[pos+25351], tapes[pos+27646], tapes[pos+29941], tapes[pos+32236], tapes[pos+34531]};
    assign tmp_shares[1727:1712]={tapes[pos+107], tapes[pos+2402], tapes[pos+4697], tapes[pos+6992], tapes[pos+9287], tapes[pos+11582], tapes[pos+13877], tapes[pos+16172], tapes[pos+18467], tapes[pos+20762], tapes[pos+23057], tapes[pos+25352], tapes[pos+27647], tapes[pos+29942], tapes[pos+32237], tapes[pos+34532]};
    assign tmp_shares[1743:1728]={tapes[pos+108], tapes[pos+2403], tapes[pos+4698], tapes[pos+6993], tapes[pos+9288], tapes[pos+11583], tapes[pos+13878], tapes[pos+16173], tapes[pos+18468], tapes[pos+20763], tapes[pos+23058], tapes[pos+25353], tapes[pos+27648], tapes[pos+29943], tapes[pos+32238], tapes[pos+34533]};
    assign tmp_shares[1759:1744]={tapes[pos+109], tapes[pos+2404], tapes[pos+4699], tapes[pos+6994], tapes[pos+9289], tapes[pos+11584], tapes[pos+13879], tapes[pos+16174], tapes[pos+18469], tapes[pos+20764], tapes[pos+23059], tapes[pos+25354], tapes[pos+27649], tapes[pos+29944], tapes[pos+32239], tapes[pos+34534]};
    assign tmp_shares[1775:1760]={tapes[pos+110], tapes[pos+2405], tapes[pos+4700], tapes[pos+6995], tapes[pos+9290], tapes[pos+11585], tapes[pos+13880], tapes[pos+16175], tapes[pos+18470], tapes[pos+20765], tapes[pos+23060], tapes[pos+25355], tapes[pos+27650], tapes[pos+29945], tapes[pos+32240], tapes[pos+34535]};
    assign tmp_shares[1791:1776]={tapes[pos+111], tapes[pos+2406], tapes[pos+4701], tapes[pos+6996], tapes[pos+9291], tapes[pos+11586], tapes[pos+13881], tapes[pos+16176], tapes[pos+18471], tapes[pos+20766], tapes[pos+23061], tapes[pos+25356], tapes[pos+27651], tapes[pos+29946], tapes[pos+32241], tapes[pos+34536]};
    assign tmp_shares[1807:1792]={tapes[pos+112], tapes[pos+2407], tapes[pos+4702], tapes[pos+6997], tapes[pos+9292], tapes[pos+11587], tapes[pos+13882], tapes[pos+16177], tapes[pos+18472], tapes[pos+20767], tapes[pos+23062], tapes[pos+25357], tapes[pos+27652], tapes[pos+29947], tapes[pos+32242], tapes[pos+34537]};
    assign tmp_shares[1823:1808]={tapes[pos+113], tapes[pos+2408], tapes[pos+4703], tapes[pos+6998], tapes[pos+9293], tapes[pos+11588], tapes[pos+13883], tapes[pos+16178], tapes[pos+18473], tapes[pos+20768], tapes[pos+23063], tapes[pos+25358], tapes[pos+27653], tapes[pos+29948], tapes[pos+32243], tapes[pos+34538]};
    assign tmp_shares[1839:1824]={tapes[pos+114], tapes[pos+2409], tapes[pos+4704], tapes[pos+6999], tapes[pos+9294], tapes[pos+11589], tapes[pos+13884], tapes[pos+16179], tapes[pos+18474], tapes[pos+20769], tapes[pos+23064], tapes[pos+25359], tapes[pos+27654], tapes[pos+29949], tapes[pos+32244], tapes[pos+34539]};
    assign tmp_shares[1855:1840]={tapes[pos+115], tapes[pos+2410], tapes[pos+4705], tapes[pos+7000], tapes[pos+9295], tapes[pos+11590], tapes[pos+13885], tapes[pos+16180], tapes[pos+18475], tapes[pos+20770], tapes[pos+23065], tapes[pos+25360], tapes[pos+27655], tapes[pos+29950], tapes[pos+32245], tapes[pos+34540]};
    assign tmp_shares[1871:1856]={tapes[pos+116], tapes[pos+2411], tapes[pos+4706], tapes[pos+7001], tapes[pos+9296], tapes[pos+11591], tapes[pos+13886], tapes[pos+16181], tapes[pos+18476], tapes[pos+20771], tapes[pos+23066], tapes[pos+25361], tapes[pos+27656], tapes[pos+29951], tapes[pos+32246], tapes[pos+34541]};
    assign tmp_shares[1887:1872]={tapes[pos+117], tapes[pos+2412], tapes[pos+4707], tapes[pos+7002], tapes[pos+9297], tapes[pos+11592], tapes[pos+13887], tapes[pos+16182], tapes[pos+18477], tapes[pos+20772], tapes[pos+23067], tapes[pos+25362], tapes[pos+27657], tapes[pos+29952], tapes[pos+32247], tapes[pos+34542]};
    assign tmp_shares[1903:1888]={tapes[pos+118], tapes[pos+2413], tapes[pos+4708], tapes[pos+7003], tapes[pos+9298], tapes[pos+11593], tapes[pos+13888], tapes[pos+16183], tapes[pos+18478], tapes[pos+20773], tapes[pos+23068], tapes[pos+25363], tapes[pos+27658], tapes[pos+29953], tapes[pos+32248], tapes[pos+34543]};
    assign tmp_shares[1919:1904]={tapes[pos+119], tapes[pos+2414], tapes[pos+4709], tapes[pos+7004], tapes[pos+9299], tapes[pos+11594], tapes[pos+13889], tapes[pos+16184], tapes[pos+18479], tapes[pos+20774], tapes[pos+23069], tapes[pos+25364], tapes[pos+27659], tapes[pos+29954], tapes[pos+32249], tapes[pos+34544]};
    assign tmp_shares[1935:1920]={tapes[pos+120], tapes[pos+2415], tapes[pos+4710], tapes[pos+7005], tapes[pos+9300], tapes[pos+11595], tapes[pos+13890], tapes[pos+16185], tapes[pos+18480], tapes[pos+20775], tapes[pos+23070], tapes[pos+25365], tapes[pos+27660], tapes[pos+29955], tapes[pos+32250], tapes[pos+34545]};
    assign tmp_shares[1951:1936]={tapes[pos+121], tapes[pos+2416], tapes[pos+4711], tapes[pos+7006], tapes[pos+9301], tapes[pos+11596], tapes[pos+13891], tapes[pos+16186], tapes[pos+18481], tapes[pos+20776], tapes[pos+23071], tapes[pos+25366], tapes[pos+27661], tapes[pos+29956], tapes[pos+32251], tapes[pos+34546]};
    assign tmp_shares[1967:1952]={tapes[pos+122], tapes[pos+2417], tapes[pos+4712], tapes[pos+7007], tapes[pos+9302], tapes[pos+11597], tapes[pos+13892], tapes[pos+16187], tapes[pos+18482], tapes[pos+20777], tapes[pos+23072], tapes[pos+25367], tapes[pos+27662], tapes[pos+29957], tapes[pos+32252], tapes[pos+34547]};
    assign tmp_shares[1983:1968]={tapes[pos+123], tapes[pos+2418], tapes[pos+4713], tapes[pos+7008], tapes[pos+9303], tapes[pos+11598], tapes[pos+13893], tapes[pos+16188], tapes[pos+18483], tapes[pos+20778], tapes[pos+23073], tapes[pos+25368], tapes[pos+27663], tapes[pos+29958], tapes[pos+32253], tapes[pos+34548]};
    assign tmp_shares[1999:1984]={tapes[pos+124], tapes[pos+2419], tapes[pos+4714], tapes[pos+7009], tapes[pos+9304], tapes[pos+11599], tapes[pos+13894], tapes[pos+16189], tapes[pos+18484], tapes[pos+20779], tapes[pos+23074], tapes[pos+25369], tapes[pos+27664], tapes[pos+29959], tapes[pos+32254], tapes[pos+34549]};
    assign tmp_shares[2015:2000]={tapes[pos+125], tapes[pos+2420], tapes[pos+4715], tapes[pos+7010], tapes[pos+9305], tapes[pos+11600], tapes[pos+13895], tapes[pos+16190], tapes[pos+18485], tapes[pos+20780], tapes[pos+23075], tapes[pos+25370], tapes[pos+27665], tapes[pos+29960], tapes[pos+32255], tapes[pos+34550]};
    assign tmp_shares[2031:2016]={tapes[pos+126], tapes[pos+2421], tapes[pos+4716], tapes[pos+7011], tapes[pos+9306], tapes[pos+11601], tapes[pos+13896], tapes[pos+16191], tapes[pos+18486], tapes[pos+20781], tapes[pos+23076], tapes[pos+25371], tapes[pos+27666], tapes[pos+29961], tapes[pos+32256], tapes[pos+34551]};
    assign tmp_shares[2047:2032]={tapes[pos+127], tapes[pos+2422], tapes[pos+4717], tapes[pos+7012], tapes[pos+9307], tapes[pos+11602], tapes[pos+13897], tapes[pos+16192], tapes[pos+18487], tapes[pos+20782], tapes[pos+23077], tapes[pos+25372], tapes[pos+27667], tapes[pos+29962], tapes[pos+32257], tapes[pos+34552]};
    assign tmp_shares[2063:2048]={tapes[pos+128], tapes[pos+2423], tapes[pos+4718], tapes[pos+7013], tapes[pos+9308], tapes[pos+11603], tapes[pos+13898], tapes[pos+16193], tapes[pos+18488], tapes[pos+20783], tapes[pos+23078], tapes[pos+25373], tapes[pos+27668], tapes[pos+29963], tapes[pos+32258], tapes[pos+34553]};
    assign tmp_shares[2079:2064]={tapes[pos+129], tapes[pos+2424], tapes[pos+4719], tapes[pos+7014], tapes[pos+9309], tapes[pos+11604], tapes[pos+13899], tapes[pos+16194], tapes[pos+18489], tapes[pos+20784], tapes[pos+23079], tapes[pos+25374], tapes[pos+27669], tapes[pos+29964], tapes[pos+32259], tapes[pos+34554]};
    assign tmp_shares[2095:2080]={tapes[pos+130], tapes[pos+2425], tapes[pos+4720], tapes[pos+7015], tapes[pos+9310], tapes[pos+11605], tapes[pos+13900], tapes[pos+16195], tapes[pos+18490], tapes[pos+20785], tapes[pos+23080], tapes[pos+25375], tapes[pos+27670], tapes[pos+29965], tapes[pos+32260], tapes[pos+34555]};
    assign tmp_shares[2111:2096]={tapes[pos+131], tapes[pos+2426], tapes[pos+4721], tapes[pos+7016], tapes[pos+9311], tapes[pos+11606], tapes[pos+13901], tapes[pos+16196], tapes[pos+18491], tapes[pos+20786], tapes[pos+23081], tapes[pos+25376], tapes[pos+27671], tapes[pos+29966], tapes[pos+32261], tapes[pos+34556]};
    assign tmp_shares[2127:2112]={tapes[pos+132], tapes[pos+2427], tapes[pos+4722], tapes[pos+7017], tapes[pos+9312], tapes[pos+11607], tapes[pos+13902], tapes[pos+16197], tapes[pos+18492], tapes[pos+20787], tapes[pos+23082], tapes[pos+25377], tapes[pos+27672], tapes[pos+29967], tapes[pos+32262], tapes[pos+34557]};
    assign tmp_shares[2143:2128]={tapes[pos+133], tapes[pos+2428], tapes[pos+4723], tapes[pos+7018], tapes[pos+9313], tapes[pos+11608], tapes[pos+13903], tapes[pos+16198], tapes[pos+18493], tapes[pos+20788], tapes[pos+23083], tapes[pos+25378], tapes[pos+27673], tapes[pos+29968], tapes[pos+32263], tapes[pos+34558]};
    assign tmp_shares[2159:2144]={tapes[pos+134], tapes[pos+2429], tapes[pos+4724], tapes[pos+7019], tapes[pos+9314], tapes[pos+11609], tapes[pos+13904], tapes[pos+16199], tapes[pos+18494], tapes[pos+20789], tapes[pos+23084], tapes[pos+25379], tapes[pos+27674], tapes[pos+29969], tapes[pos+32264], tapes[pos+34559]};
    assign tmp_shares[2175:2160]={tapes[pos+135], tapes[pos+2430], tapes[pos+4725], tapes[pos+7020], tapes[pos+9315], tapes[pos+11610], tapes[pos+13905], tapes[pos+16200], tapes[pos+18495], tapes[pos+20790], tapes[pos+23085], tapes[pos+25380], tapes[pos+27675], tapes[pos+29970], tapes[pos+32265], tapes[pos+34560]};
    assign tmp_shares[2191:2176]={tapes[pos+136], tapes[pos+2431], tapes[pos+4726], tapes[pos+7021], tapes[pos+9316], tapes[pos+11611], tapes[pos+13906], tapes[pos+16201], tapes[pos+18496], tapes[pos+20791], tapes[pos+23086], tapes[pos+25381], tapes[pos+27676], tapes[pos+29971], tapes[pos+32266], tapes[pos+34561]};
    assign tmp_shares[2207:2192]={tapes[pos+137], tapes[pos+2432], tapes[pos+4727], tapes[pos+7022], tapes[pos+9317], tapes[pos+11612], tapes[pos+13907], tapes[pos+16202], tapes[pos+18497], tapes[pos+20792], tapes[pos+23087], tapes[pos+25382], tapes[pos+27677], tapes[pos+29972], tapes[pos+32267], tapes[pos+34562]};
    assign tmp_shares[2223:2208]={tapes[pos+138], tapes[pos+2433], tapes[pos+4728], tapes[pos+7023], tapes[pos+9318], tapes[pos+11613], tapes[pos+13908], tapes[pos+16203], tapes[pos+18498], tapes[pos+20793], tapes[pos+23088], tapes[pos+25383], tapes[pos+27678], tapes[pos+29973], tapes[pos+32268], tapes[pos+34563]};
    assign tmp_shares[2239:2224]={tapes[pos+139], tapes[pos+2434], tapes[pos+4729], tapes[pos+7024], tapes[pos+9319], tapes[pos+11614], tapes[pos+13909], tapes[pos+16204], tapes[pos+18499], tapes[pos+20794], tapes[pos+23089], tapes[pos+25384], tapes[pos+27679], tapes[pos+29974], tapes[pos+32269], tapes[pos+34564]};
    assign tmp_shares[2255:2240]={tapes[pos+140], tapes[pos+2435], tapes[pos+4730], tapes[pos+7025], tapes[pos+9320], tapes[pos+11615], tapes[pos+13910], tapes[pos+16205], tapes[pos+18500], tapes[pos+20795], tapes[pos+23090], tapes[pos+25385], tapes[pos+27680], tapes[pos+29975], tapes[pos+32270], tapes[pos+34565]};
    assign tmp_shares[2271:2256]={tapes[pos+141], tapes[pos+2436], tapes[pos+4731], tapes[pos+7026], tapes[pos+9321], tapes[pos+11616], tapes[pos+13911], tapes[pos+16206], tapes[pos+18501], tapes[pos+20796], tapes[pos+23091], tapes[pos+25386], tapes[pos+27681], tapes[pos+29976], tapes[pos+32271], tapes[pos+34566]};
    assign tmp_shares[2287:2272]={tapes[pos+142], tapes[pos+2437], tapes[pos+4732], tapes[pos+7027], tapes[pos+9322], tapes[pos+11617], tapes[pos+13912], tapes[pos+16207], tapes[pos+18502], tapes[pos+20797], tapes[pos+23092], tapes[pos+25387], tapes[pos+27682], tapes[pos+29977], tapes[pos+32272], tapes[pos+34567]};
    assign tmp_shares[2303:2288]={tapes[pos+143], tapes[pos+2438], tapes[pos+4733], tapes[pos+7028], tapes[pos+9323], tapes[pos+11618], tapes[pos+13913], tapes[pos+16208], tapes[pos+18503], tapes[pos+20798], tapes[pos+23093], tapes[pos+25388], tapes[pos+27683], tapes[pos+29978], tapes[pos+32273], tapes[pos+34568]};
    assign tmp_shares[2319:2304]={tapes[pos+144], tapes[pos+2439], tapes[pos+4734], tapes[pos+7029], tapes[pos+9324], tapes[pos+11619], tapes[pos+13914], tapes[pos+16209], tapes[pos+18504], tapes[pos+20799], tapes[pos+23094], tapes[pos+25389], tapes[pos+27684], tapes[pos+29979], tapes[pos+32274], tapes[pos+34569]};
    assign tmp_shares[2335:2320]={tapes[pos+145], tapes[pos+2440], tapes[pos+4735], tapes[pos+7030], tapes[pos+9325], tapes[pos+11620], tapes[pos+13915], tapes[pos+16210], tapes[pos+18505], tapes[pos+20800], tapes[pos+23095], tapes[pos+25390], tapes[pos+27685], tapes[pos+29980], tapes[pos+32275], tapes[pos+34570]};
    assign tmp_shares[2351:2336]={tapes[pos+146], tapes[pos+2441], tapes[pos+4736], tapes[pos+7031], tapes[pos+9326], tapes[pos+11621], tapes[pos+13916], tapes[pos+16211], tapes[pos+18506], tapes[pos+20801], tapes[pos+23096], tapes[pos+25391], tapes[pos+27686], tapes[pos+29981], tapes[pos+32276], tapes[pos+34571]};
    assign tmp_shares[2367:2352]={tapes[pos+147], tapes[pos+2442], tapes[pos+4737], tapes[pos+7032], tapes[pos+9327], tapes[pos+11622], tapes[pos+13917], tapes[pos+16212], tapes[pos+18507], tapes[pos+20802], tapes[pos+23097], tapes[pos+25392], tapes[pos+27687], tapes[pos+29982], tapes[pos+32277], tapes[pos+34572]};
    assign tmp_shares[2383:2368]={tapes[pos+148], tapes[pos+2443], tapes[pos+4738], tapes[pos+7033], tapes[pos+9328], tapes[pos+11623], tapes[pos+13918], tapes[pos+16213], tapes[pos+18508], tapes[pos+20803], tapes[pos+23098], tapes[pos+25393], tapes[pos+27688], tapes[pos+29983], tapes[pos+32278], tapes[pos+34573]};
    assign tmp_shares[2399:2384]={tapes[pos+149], tapes[pos+2444], tapes[pos+4739], tapes[pos+7034], tapes[pos+9329], tapes[pos+11624], tapes[pos+13919], tapes[pos+16214], tapes[pos+18509], tapes[pos+20804], tapes[pos+23099], tapes[pos+25394], tapes[pos+27689], tapes[pos+29984], tapes[pos+32279], tapes[pos+34574]};
    assign tmp_shares[2415:2400]={tapes[pos+150], tapes[pos+2445], tapes[pos+4740], tapes[pos+7035], tapes[pos+9330], tapes[pos+11625], tapes[pos+13920], tapes[pos+16215], tapes[pos+18510], tapes[pos+20805], tapes[pos+23100], tapes[pos+25395], tapes[pos+27690], tapes[pos+29985], tapes[pos+32280], tapes[pos+34575]};
    assign tmp_shares[2431:2416]={tapes[pos+151], tapes[pos+2446], tapes[pos+4741], tapes[pos+7036], tapes[pos+9331], tapes[pos+11626], tapes[pos+13921], tapes[pos+16216], tapes[pos+18511], tapes[pos+20806], tapes[pos+23101], tapes[pos+25396], tapes[pos+27691], tapes[pos+29986], tapes[pos+32281], tapes[pos+34576]};
    assign tmp_shares[2447:2432]={tapes[pos+152], tapes[pos+2447], tapes[pos+4742], tapes[pos+7037], tapes[pos+9332], tapes[pos+11627], tapes[pos+13922], tapes[pos+16217], tapes[pos+18512], tapes[pos+20807], tapes[pos+23102], tapes[pos+25397], tapes[pos+27692], tapes[pos+29987], tapes[pos+32282], tapes[pos+34577]};
    assign tmp_shares[2463:2448]={tapes[pos+153], tapes[pos+2448], tapes[pos+4743], tapes[pos+7038], tapes[pos+9333], tapes[pos+11628], tapes[pos+13923], tapes[pos+16218], tapes[pos+18513], tapes[pos+20808], tapes[pos+23103], tapes[pos+25398], tapes[pos+27693], tapes[pos+29988], tapes[pos+32283], tapes[pos+34578]};
    assign tmp_shares[2479:2464]={tapes[pos+154], tapes[pos+2449], tapes[pos+4744], tapes[pos+7039], tapes[pos+9334], tapes[pos+11629], tapes[pos+13924], tapes[pos+16219], tapes[pos+18514], tapes[pos+20809], tapes[pos+23104], tapes[pos+25399], tapes[pos+27694], tapes[pos+29989], tapes[pos+32284], tapes[pos+34579]};
    assign tmp_shares[2495:2480]={tapes[pos+155], tapes[pos+2450], tapes[pos+4745], tapes[pos+7040], tapes[pos+9335], tapes[pos+11630], tapes[pos+13925], tapes[pos+16220], tapes[pos+18515], tapes[pos+20810], tapes[pos+23105], tapes[pos+25400], tapes[pos+27695], tapes[pos+29990], tapes[pos+32285], tapes[pos+34580]};
    assign tmp_shares[2511:2496]={tapes[pos+156], tapes[pos+2451], tapes[pos+4746], tapes[pos+7041], tapes[pos+9336], tapes[pos+11631], tapes[pos+13926], tapes[pos+16221], tapes[pos+18516], tapes[pos+20811], tapes[pos+23106], tapes[pos+25401], tapes[pos+27696], tapes[pos+29991], tapes[pos+32286], tapes[pos+34581]};
    assign tmp_shares[2527:2512]={tapes[pos+157], tapes[pos+2452], tapes[pos+4747], tapes[pos+7042], tapes[pos+9337], tapes[pos+11632], tapes[pos+13927], tapes[pos+16222], tapes[pos+18517], tapes[pos+20812], tapes[pos+23107], tapes[pos+25402], tapes[pos+27697], tapes[pos+29992], tapes[pos+32287], tapes[pos+34582]};
    assign tmp_shares[2543:2528]={tapes[pos+158], tapes[pos+2453], tapes[pos+4748], tapes[pos+7043], tapes[pos+9338], tapes[pos+11633], tapes[pos+13928], tapes[pos+16223], tapes[pos+18518], tapes[pos+20813], tapes[pos+23108], tapes[pos+25403], tapes[pos+27698], tapes[pos+29993], tapes[pos+32288], tapes[pos+34583]};
    assign tmp_shares[2559:2544]={tapes[pos+159], tapes[pos+2454], tapes[pos+4749], tapes[pos+7044], tapes[pos+9339], tapes[pos+11634], tapes[pos+13929], tapes[pos+16224], tapes[pos+18519], tapes[pos+20814], tapes[pos+23109], tapes[pos+25404], tapes[pos+27699], tapes[pos+29994], tapes[pos+32289], tapes[pos+34584]};
    assign tmp_shares[2575:2560]={tapes[pos+160], tapes[pos+2455], tapes[pos+4750], tapes[pos+7045], tapes[pos+9340], tapes[pos+11635], tapes[pos+13930], tapes[pos+16225], tapes[pos+18520], tapes[pos+20815], tapes[pos+23110], tapes[pos+25405], tapes[pos+27700], tapes[pos+29995], tapes[pos+32290], tapes[pos+34585]};
    assign tmp_shares[2591:2576]={tapes[pos+161], tapes[pos+2456], tapes[pos+4751], tapes[pos+7046], tapes[pos+9341], tapes[pos+11636], tapes[pos+13931], tapes[pos+16226], tapes[pos+18521], tapes[pos+20816], tapes[pos+23111], tapes[pos+25406], tapes[pos+27701], tapes[pos+29996], tapes[pos+32291], tapes[pos+34586]};
    assign tmp_shares[2607:2592]={tapes[pos+162], tapes[pos+2457], tapes[pos+4752], tapes[pos+7047], tapes[pos+9342], tapes[pos+11637], tapes[pos+13932], tapes[pos+16227], tapes[pos+18522], tapes[pos+20817], tapes[pos+23112], tapes[pos+25407], tapes[pos+27702], tapes[pos+29997], tapes[pos+32292], tapes[pos+34587]};
    assign tmp_shares[2623:2608]={tapes[pos+163], tapes[pos+2458], tapes[pos+4753], tapes[pos+7048], tapes[pos+9343], tapes[pos+11638], tapes[pos+13933], tapes[pos+16228], tapes[pos+18523], tapes[pos+20818], tapes[pos+23113], tapes[pos+25408], tapes[pos+27703], tapes[pos+29998], tapes[pos+32293], tapes[pos+34588]};
    assign tmp_shares[2639:2624]={tapes[pos+164], tapes[pos+2459], tapes[pos+4754], tapes[pos+7049], tapes[pos+9344], tapes[pos+11639], tapes[pos+13934], tapes[pos+16229], tapes[pos+18524], tapes[pos+20819], tapes[pos+23114], tapes[pos+25409], tapes[pos+27704], tapes[pos+29999], tapes[pos+32294], tapes[pos+34589]};
    assign tmp_shares[2655:2640]={tapes[pos+165], tapes[pos+2460], tapes[pos+4755], tapes[pos+7050], tapes[pos+9345], tapes[pos+11640], tapes[pos+13935], tapes[pos+16230], tapes[pos+18525], tapes[pos+20820], tapes[pos+23115], tapes[pos+25410], tapes[pos+27705], tapes[pos+30000], tapes[pos+32295], tapes[pos+34590]};
    assign tmp_shares[2671:2656]={tapes[pos+166], tapes[pos+2461], tapes[pos+4756], tapes[pos+7051], tapes[pos+9346], tapes[pos+11641], tapes[pos+13936], tapes[pos+16231], tapes[pos+18526], tapes[pos+20821], tapes[pos+23116], tapes[pos+25411], tapes[pos+27706], tapes[pos+30001], tapes[pos+32296], tapes[pos+34591]};
    assign tmp_shares[2687:2672]={tapes[pos+167], tapes[pos+2462], tapes[pos+4757], tapes[pos+7052], tapes[pos+9347], tapes[pos+11642], tapes[pos+13937], tapes[pos+16232], tapes[pos+18527], tapes[pos+20822], tapes[pos+23117], tapes[pos+25412], tapes[pos+27707], tapes[pos+30002], tapes[pos+32297], tapes[pos+34592]};
    assign tmp_shares[2703:2688]={tapes[pos+168], tapes[pos+2463], tapes[pos+4758], tapes[pos+7053], tapes[pos+9348], tapes[pos+11643], tapes[pos+13938], tapes[pos+16233], tapes[pos+18528], tapes[pos+20823], tapes[pos+23118], tapes[pos+25413], tapes[pos+27708], tapes[pos+30003], tapes[pos+32298], tapes[pos+34593]};
    assign tmp_shares[2719:2704]={tapes[pos+169], tapes[pos+2464], tapes[pos+4759], tapes[pos+7054], tapes[pos+9349], tapes[pos+11644], tapes[pos+13939], tapes[pos+16234], tapes[pos+18529], tapes[pos+20824], tapes[pos+23119], tapes[pos+25414], tapes[pos+27709], tapes[pos+30004], tapes[pos+32299], tapes[pos+34594]};
    assign tmp_shares[2735:2720]={tapes[pos+170], tapes[pos+2465], tapes[pos+4760], tapes[pos+7055], tapes[pos+9350], tapes[pos+11645], tapes[pos+13940], tapes[pos+16235], tapes[pos+18530], tapes[pos+20825], tapes[pos+23120], tapes[pos+25415], tapes[pos+27710], tapes[pos+30005], tapes[pos+32300], tapes[pos+34595]};
    assign tmp_shares[2751:2736]={tapes[pos+171], tapes[pos+2466], tapes[pos+4761], tapes[pos+7056], tapes[pos+9351], tapes[pos+11646], tapes[pos+13941], tapes[pos+16236], tapes[pos+18531], tapes[pos+20826], tapes[pos+23121], tapes[pos+25416], tapes[pos+27711], tapes[pos+30006], tapes[pos+32301], tapes[pos+34596]};
    assign tmp_shares[2767:2752]={tapes[pos+172], tapes[pos+2467], tapes[pos+4762], tapes[pos+7057], tapes[pos+9352], tapes[pos+11647], tapes[pos+13942], tapes[pos+16237], tapes[pos+18532], tapes[pos+20827], tapes[pos+23122], tapes[pos+25417], tapes[pos+27712], tapes[pos+30007], tapes[pos+32302], tapes[pos+34597]};
    assign tmp_shares[2783:2768]={tapes[pos+173], tapes[pos+2468], tapes[pos+4763], tapes[pos+7058], tapes[pos+9353], tapes[pos+11648], tapes[pos+13943], tapes[pos+16238], tapes[pos+18533], tapes[pos+20828], tapes[pos+23123], tapes[pos+25418], tapes[pos+27713], tapes[pos+30008], tapes[pos+32303], tapes[pos+34598]};
    assign tmp_shares[2799:2784]={tapes[pos+174], tapes[pos+2469], tapes[pos+4764], tapes[pos+7059], tapes[pos+9354], tapes[pos+11649], tapes[pos+13944], tapes[pos+16239], tapes[pos+18534], tapes[pos+20829], tapes[pos+23124], tapes[pos+25419], tapes[pos+27714], tapes[pos+30009], tapes[pos+32304], tapes[pos+34599]};
    assign tmp_shares[2815:2800]={tapes[pos+175], tapes[pos+2470], tapes[pos+4765], tapes[pos+7060], tapes[pos+9355], tapes[pos+11650], tapes[pos+13945], tapes[pos+16240], tapes[pos+18535], tapes[pos+20830], tapes[pos+23125], tapes[pos+25420], tapes[pos+27715], tapes[pos+30010], tapes[pos+32305], tapes[pos+34600]};
    assign tmp_shares[2831:2816]={tapes[pos+176], tapes[pos+2471], tapes[pos+4766], tapes[pos+7061], tapes[pos+9356], tapes[pos+11651], tapes[pos+13946], tapes[pos+16241], tapes[pos+18536], tapes[pos+20831], tapes[pos+23126], tapes[pos+25421], tapes[pos+27716], tapes[pos+30011], tapes[pos+32306], tapes[pos+34601]};
    assign tmp_shares[2847:2832]={tapes[pos+177], tapes[pos+2472], tapes[pos+4767], tapes[pos+7062], tapes[pos+9357], tapes[pos+11652], tapes[pos+13947], tapes[pos+16242], tapes[pos+18537], tapes[pos+20832], tapes[pos+23127], tapes[pos+25422], tapes[pos+27717], tapes[pos+30012], tapes[pos+32307], tapes[pos+34602]};
    assign tmp_shares[2863:2848]={tapes[pos+178], tapes[pos+2473], tapes[pos+4768], tapes[pos+7063], tapes[pos+9358], tapes[pos+11653], tapes[pos+13948], tapes[pos+16243], tapes[pos+18538], tapes[pos+20833], tapes[pos+23128], tapes[pos+25423], tapes[pos+27718], tapes[pos+30013], tapes[pos+32308], tapes[pos+34603]};
    assign tmp_shares[2879:2864]={tapes[pos+179], tapes[pos+2474], tapes[pos+4769], tapes[pos+7064], tapes[pos+9359], tapes[pos+11654], tapes[pos+13949], tapes[pos+16244], tapes[pos+18539], tapes[pos+20834], tapes[pos+23129], tapes[pos+25424], tapes[pos+27719], tapes[pos+30014], tapes[pos+32309], tapes[pos+34604]};
    assign tmp_shares[2895:2880]={tapes[pos+180], tapes[pos+2475], tapes[pos+4770], tapes[pos+7065], tapes[pos+9360], tapes[pos+11655], tapes[pos+13950], tapes[pos+16245], tapes[pos+18540], tapes[pos+20835], tapes[pos+23130], tapes[pos+25425], tapes[pos+27720], tapes[pos+30015], tapes[pos+32310], tapes[pos+34605]};
    assign tmp_shares[2911:2896]={tapes[pos+181], tapes[pos+2476], tapes[pos+4771], tapes[pos+7066], tapes[pos+9361], tapes[pos+11656], tapes[pos+13951], tapes[pos+16246], tapes[pos+18541], tapes[pos+20836], tapes[pos+23131], tapes[pos+25426], tapes[pos+27721], tapes[pos+30016], tapes[pos+32311], tapes[pos+34606]};
    assign tmp_shares[2927:2912]={tapes[pos+182], tapes[pos+2477], tapes[pos+4772], tapes[pos+7067], tapes[pos+9362], tapes[pos+11657], tapes[pos+13952], tapes[pos+16247], tapes[pos+18542], tapes[pos+20837], tapes[pos+23132], tapes[pos+25427], tapes[pos+27722], tapes[pos+30017], tapes[pos+32312], tapes[pos+34607]};
    assign tmp_shares[2943:2928]={tapes[pos+183], tapes[pos+2478], tapes[pos+4773], tapes[pos+7068], tapes[pos+9363], tapes[pos+11658], tapes[pos+13953], tapes[pos+16248], tapes[pos+18543], tapes[pos+20838], tapes[pos+23133], tapes[pos+25428], tapes[pos+27723], tapes[pos+30018], tapes[pos+32313], tapes[pos+34608]};
    assign tmp_shares[2959:2944]={tapes[pos+184], tapes[pos+2479], tapes[pos+4774], tapes[pos+7069], tapes[pos+9364], tapes[pos+11659], tapes[pos+13954], tapes[pos+16249], tapes[pos+18544], tapes[pos+20839], tapes[pos+23134], tapes[pos+25429], tapes[pos+27724], tapes[pos+30019], tapes[pos+32314], tapes[pos+34609]};
    assign tmp_shares[2975:2960]={tapes[pos+185], tapes[pos+2480], tapes[pos+4775], tapes[pos+7070], tapes[pos+9365], tapes[pos+11660], tapes[pos+13955], tapes[pos+16250], tapes[pos+18545], tapes[pos+20840], tapes[pos+23135], tapes[pos+25430], tapes[pos+27725], tapes[pos+30020], tapes[pos+32315], tapes[pos+34610]};
    assign tmp_shares[2991:2976]={tapes[pos+186], tapes[pos+2481], tapes[pos+4776], tapes[pos+7071], tapes[pos+9366], tapes[pos+11661], tapes[pos+13956], tapes[pos+16251], tapes[pos+18546], tapes[pos+20841], tapes[pos+23136], tapes[pos+25431], tapes[pos+27726], tapes[pos+30021], tapes[pos+32316], tapes[pos+34611]};
    assign tmp_shares[3007:2992]={tapes[pos+187], tapes[pos+2482], tapes[pos+4777], tapes[pos+7072], tapes[pos+9367], tapes[pos+11662], tapes[pos+13957], tapes[pos+16252], tapes[pos+18547], tapes[pos+20842], tapes[pos+23137], tapes[pos+25432], tapes[pos+27727], tapes[pos+30022], tapes[pos+32317], tapes[pos+34612]};
    assign tmp_shares[3023:3008]={tapes[pos+188], tapes[pos+2483], tapes[pos+4778], tapes[pos+7073], tapes[pos+9368], tapes[pos+11663], tapes[pos+13958], tapes[pos+16253], tapes[pos+18548], tapes[pos+20843], tapes[pos+23138], tapes[pos+25433], tapes[pos+27728], tapes[pos+30023], tapes[pos+32318], tapes[pos+34613]};
    assign tmp_shares[3039:3024]={tapes[pos+189], tapes[pos+2484], tapes[pos+4779], tapes[pos+7074], tapes[pos+9369], tapes[pos+11664], tapes[pos+13959], tapes[pos+16254], tapes[pos+18549], tapes[pos+20844], tapes[pos+23139], tapes[pos+25434], tapes[pos+27729], tapes[pos+30024], tapes[pos+32319], tapes[pos+34614]};
    assign tmp_shares[3055:3040]={tapes[pos+190], tapes[pos+2485], tapes[pos+4780], tapes[pos+7075], tapes[pos+9370], tapes[pos+11665], tapes[pos+13960], tapes[pos+16255], tapes[pos+18550], tapes[pos+20845], tapes[pos+23140], tapes[pos+25435], tapes[pos+27730], tapes[pos+30025], tapes[pos+32320], tapes[pos+34615]};
    assign tmp_shares[3071:3056]={tapes[pos+191], tapes[pos+2486], tapes[pos+4781], tapes[pos+7076], tapes[pos+9371], tapes[pos+11666], tapes[pos+13961], tapes[pos+16256], tapes[pos+18551], tapes[pos+20846], tapes[pos+23141], tapes[pos+25436], tapes[pos+27731], tapes[pos+30026], tapes[pos+32321], tapes[pos+34616]};
    assign tmp_shares[3087:3072]={tapes[pos+192], tapes[pos+2487], tapes[pos+4782], tapes[pos+7077], tapes[pos+9372], tapes[pos+11667], tapes[pos+13962], tapes[pos+16257], tapes[pos+18552], tapes[pos+20847], tapes[pos+23142], tapes[pos+25437], tapes[pos+27732], tapes[pos+30027], tapes[pos+32322], tapes[pos+34617]};
    assign tmp_shares[3103:3088]={tapes[pos+193], tapes[pos+2488], tapes[pos+4783], tapes[pos+7078], tapes[pos+9373], tapes[pos+11668], tapes[pos+13963], tapes[pos+16258], tapes[pos+18553], tapes[pos+20848], tapes[pos+23143], tapes[pos+25438], tapes[pos+27733], tapes[pos+30028], tapes[pos+32323], tapes[pos+34618]};
    assign tmp_shares[3119:3104]={tapes[pos+194], tapes[pos+2489], tapes[pos+4784], tapes[pos+7079], tapes[pos+9374], tapes[pos+11669], tapes[pos+13964], tapes[pos+16259], tapes[pos+18554], tapes[pos+20849], tapes[pos+23144], tapes[pos+25439], tapes[pos+27734], tapes[pos+30029], tapes[pos+32324], tapes[pos+34619]};
    assign tmp_shares[3135:3120]={tapes[pos+195], tapes[pos+2490], tapes[pos+4785], tapes[pos+7080], tapes[pos+9375], tapes[pos+11670], tapes[pos+13965], tapes[pos+16260], tapes[pos+18555], tapes[pos+20850], tapes[pos+23145], tapes[pos+25440], tapes[pos+27735], tapes[pos+30030], tapes[pos+32325], tapes[pos+34620]};
    assign tmp_shares[3151:3136]={tapes[pos+196], tapes[pos+2491], tapes[pos+4786], tapes[pos+7081], tapes[pos+9376], tapes[pos+11671], tapes[pos+13966], tapes[pos+16261], tapes[pos+18556], tapes[pos+20851], tapes[pos+23146], tapes[pos+25441], tapes[pos+27736], tapes[pos+30031], tapes[pos+32326], tapes[pos+34621]};
    assign tmp_shares[3167:3152]={tapes[pos+197], tapes[pos+2492], tapes[pos+4787], tapes[pos+7082], tapes[pos+9377], tapes[pos+11672], tapes[pos+13967], tapes[pos+16262], tapes[pos+18557], tapes[pos+20852], tapes[pos+23147], tapes[pos+25442], tapes[pos+27737], tapes[pos+30032], tapes[pos+32327], tapes[pos+34622]};
    assign tmp_shares[3183:3168]={tapes[pos+198], tapes[pos+2493], tapes[pos+4788], tapes[pos+7083], tapes[pos+9378], tapes[pos+11673], tapes[pos+13968], tapes[pos+16263], tapes[pos+18558], tapes[pos+20853], tapes[pos+23148], tapes[pos+25443], tapes[pos+27738], tapes[pos+30033], tapes[pos+32328], tapes[pos+34623]};
    assign tmp_shares[3199:3184]={tapes[pos+199], tapes[pos+2494], tapes[pos+4789], tapes[pos+7084], tapes[pos+9379], tapes[pos+11674], tapes[pos+13969], tapes[pos+16264], tapes[pos+18559], tapes[pos+20854], tapes[pos+23149], tapes[pos+25444], tapes[pos+27739], tapes[pos+30034], tapes[pos+32329], tapes[pos+34624]};
    assign tmp_shares[3215:3200]={tapes[pos+200], tapes[pos+2495], tapes[pos+4790], tapes[pos+7085], tapes[pos+9380], tapes[pos+11675], tapes[pos+13970], tapes[pos+16265], tapes[pos+18560], tapes[pos+20855], tapes[pos+23150], tapes[pos+25445], tapes[pos+27740], tapes[pos+30035], tapes[pos+32330], tapes[pos+34625]};
    assign tmp_shares[3231:3216]={tapes[pos+201], tapes[pos+2496], tapes[pos+4791], tapes[pos+7086], tapes[pos+9381], tapes[pos+11676], tapes[pos+13971], tapes[pos+16266], tapes[pos+18561], tapes[pos+20856], tapes[pos+23151], tapes[pos+25446], tapes[pos+27741], tapes[pos+30036], tapes[pos+32331], tapes[pos+34626]};
    assign tmp_shares[3247:3232]={tapes[pos+202], tapes[pos+2497], tapes[pos+4792], tapes[pos+7087], tapes[pos+9382], tapes[pos+11677], tapes[pos+13972], tapes[pos+16267], tapes[pos+18562], tapes[pos+20857], tapes[pos+23152], tapes[pos+25447], tapes[pos+27742], tapes[pos+30037], tapes[pos+32332], tapes[pos+34627]};
    assign tmp_shares[3263:3248]={tapes[pos+203], tapes[pos+2498], tapes[pos+4793], tapes[pos+7088], tapes[pos+9383], tapes[pos+11678], tapes[pos+13973], tapes[pos+16268], tapes[pos+18563], tapes[pos+20858], tapes[pos+23153], tapes[pos+25448], tapes[pos+27743], tapes[pos+30038], tapes[pos+32333], tapes[pos+34628]};
    assign tmp_shares[3279:3264]={tapes[pos+204], tapes[pos+2499], tapes[pos+4794], tapes[pos+7089], tapes[pos+9384], tapes[pos+11679], tapes[pos+13974], tapes[pos+16269], tapes[pos+18564], tapes[pos+20859], tapes[pos+23154], tapes[pos+25449], tapes[pos+27744], tapes[pos+30039], tapes[pos+32334], tapes[pos+34629]};
    assign tmp_shares[3295:3280]={tapes[pos+205], tapes[pos+2500], tapes[pos+4795], tapes[pos+7090], tapes[pos+9385], tapes[pos+11680], tapes[pos+13975], tapes[pos+16270], tapes[pos+18565], tapes[pos+20860], tapes[pos+23155], tapes[pos+25450], tapes[pos+27745], tapes[pos+30040], tapes[pos+32335], tapes[pos+34630]};
    assign tmp_shares[3311:3296]={tapes[pos+206], tapes[pos+2501], tapes[pos+4796], tapes[pos+7091], tapes[pos+9386], tapes[pos+11681], tapes[pos+13976], tapes[pos+16271], tapes[pos+18566], tapes[pos+20861], tapes[pos+23156], tapes[pos+25451], tapes[pos+27746], tapes[pos+30041], tapes[pos+32336], tapes[pos+34631]};
    assign tmp_shares[3327:3312]={tapes[pos+207], tapes[pos+2502], tapes[pos+4797], tapes[pos+7092], tapes[pos+9387], tapes[pos+11682], tapes[pos+13977], tapes[pos+16272], tapes[pos+18567], tapes[pos+20862], tapes[pos+23157], tapes[pos+25452], tapes[pos+27747], tapes[pos+30042], tapes[pos+32337], tapes[pos+34632]};
    assign tmp_shares[3343:3328]={tapes[pos+208], tapes[pos+2503], tapes[pos+4798], tapes[pos+7093], tapes[pos+9388], tapes[pos+11683], tapes[pos+13978], tapes[pos+16273], tapes[pos+18568], tapes[pos+20863], tapes[pos+23158], tapes[pos+25453], tapes[pos+27748], tapes[pos+30043], tapes[pos+32338], tapes[pos+34633]};
    assign tmp_shares[3359:3344]={tapes[pos+209], tapes[pos+2504], tapes[pos+4799], tapes[pos+7094], tapes[pos+9389], tapes[pos+11684], tapes[pos+13979], tapes[pos+16274], tapes[pos+18569], tapes[pos+20864], tapes[pos+23159], tapes[pos+25454], tapes[pos+27749], tapes[pos+30044], tapes[pos+32339], tapes[pos+34634]};
    assign tmp_shares[3375:3360]={tapes[pos+210], tapes[pos+2505], tapes[pos+4800], tapes[pos+7095], tapes[pos+9390], tapes[pos+11685], tapes[pos+13980], tapes[pos+16275], tapes[pos+18570], tapes[pos+20865], tapes[pos+23160], tapes[pos+25455], tapes[pos+27750], tapes[pos+30045], tapes[pos+32340], tapes[pos+34635]};
    assign tmp_shares[3391:3376]={tapes[pos+211], tapes[pos+2506], tapes[pos+4801], tapes[pos+7096], tapes[pos+9391], tapes[pos+11686], tapes[pos+13981], tapes[pos+16276], tapes[pos+18571], tapes[pos+20866], tapes[pos+23161], tapes[pos+25456], tapes[pos+27751], tapes[pos+30046], tapes[pos+32341], tapes[pos+34636]};
    assign tmp_shares[3407:3392]={tapes[pos+212], tapes[pos+2507], tapes[pos+4802], tapes[pos+7097], tapes[pos+9392], tapes[pos+11687], tapes[pos+13982], tapes[pos+16277], tapes[pos+18572], tapes[pos+20867], tapes[pos+23162], tapes[pos+25457], tapes[pos+27752], tapes[pos+30047], tapes[pos+32342], tapes[pos+34637]};
    assign tmp_shares[3423:3408]={tapes[pos+213], tapes[pos+2508], tapes[pos+4803], tapes[pos+7098], tapes[pos+9393], tapes[pos+11688], tapes[pos+13983], tapes[pos+16278], tapes[pos+18573], tapes[pos+20868], tapes[pos+23163], tapes[pos+25458], tapes[pos+27753], tapes[pos+30048], tapes[pos+32343], tapes[pos+34638]};
    assign tmp_shares[3439:3424]={tapes[pos+214], tapes[pos+2509], tapes[pos+4804], tapes[pos+7099], tapes[pos+9394], tapes[pos+11689], tapes[pos+13984], tapes[pos+16279], tapes[pos+18574], tapes[pos+20869], tapes[pos+23164], tapes[pos+25459], tapes[pos+27754], tapes[pos+30049], tapes[pos+32344], tapes[pos+34639]};
    assign tmp_shares[3455:3440]={tapes[pos+215], tapes[pos+2510], tapes[pos+4805], tapes[pos+7100], tapes[pos+9395], tapes[pos+11690], tapes[pos+13985], tapes[pos+16280], tapes[pos+18575], tapes[pos+20870], tapes[pos+23165], tapes[pos+25460], tapes[pos+27755], tapes[pos+30050], tapes[pos+32345], tapes[pos+34640]};
    assign tmp_shares[3471:3456]={tapes[pos+216], tapes[pos+2511], tapes[pos+4806], tapes[pos+7101], tapes[pos+9396], tapes[pos+11691], tapes[pos+13986], tapes[pos+16281], tapes[pos+18576], tapes[pos+20871], tapes[pos+23166], tapes[pos+25461], tapes[pos+27756], tapes[pos+30051], tapes[pos+32346], tapes[pos+34641]};
    assign tmp_shares[3487:3472]={tapes[pos+217], tapes[pos+2512], tapes[pos+4807], tapes[pos+7102], tapes[pos+9397], tapes[pos+11692], tapes[pos+13987], tapes[pos+16282], tapes[pos+18577], tapes[pos+20872], tapes[pos+23167], tapes[pos+25462], tapes[pos+27757], tapes[pos+30052], tapes[pos+32347], tapes[pos+34642]};
    assign tmp_shares[3503:3488]={tapes[pos+218], tapes[pos+2513], tapes[pos+4808], tapes[pos+7103], tapes[pos+9398], tapes[pos+11693], tapes[pos+13988], tapes[pos+16283], tapes[pos+18578], tapes[pos+20873], tapes[pos+23168], tapes[pos+25463], tapes[pos+27758], tapes[pos+30053], tapes[pos+32348], tapes[pos+34643]};
    assign tmp_shares[3519:3504]={tapes[pos+219], tapes[pos+2514], tapes[pos+4809], tapes[pos+7104], tapes[pos+9399], tapes[pos+11694], tapes[pos+13989], tapes[pos+16284], tapes[pos+18579], tapes[pos+20874], tapes[pos+23169], tapes[pos+25464], tapes[pos+27759], tapes[pos+30054], tapes[pos+32349], tapes[pos+34644]};
    assign tmp_shares[3535:3520]={tapes[pos+220], tapes[pos+2515], tapes[pos+4810], tapes[pos+7105], tapes[pos+9400], tapes[pos+11695], tapes[pos+13990], tapes[pos+16285], tapes[pos+18580], tapes[pos+20875], tapes[pos+23170], tapes[pos+25465], tapes[pos+27760], tapes[pos+30055], tapes[pos+32350], tapes[pos+34645]};
    assign tmp_shares[3551:3536]={tapes[pos+221], tapes[pos+2516], tapes[pos+4811], tapes[pos+7106], tapes[pos+9401], tapes[pos+11696], tapes[pos+13991], tapes[pos+16286], tapes[pos+18581], tapes[pos+20876], tapes[pos+23171], tapes[pos+25466], tapes[pos+27761], tapes[pos+30056], tapes[pos+32351], tapes[pos+34646]};
    assign tmp_shares[3567:3552]={tapes[pos+222], tapes[pos+2517], tapes[pos+4812], tapes[pos+7107], tapes[pos+9402], tapes[pos+11697], tapes[pos+13992], tapes[pos+16287], tapes[pos+18582], tapes[pos+20877], tapes[pos+23172], tapes[pos+25467], tapes[pos+27762], tapes[pos+30057], tapes[pos+32352], tapes[pos+34647]};
    assign tmp_shares[3583:3568]={tapes[pos+223], tapes[pos+2518], tapes[pos+4813], tapes[pos+7108], tapes[pos+9403], tapes[pos+11698], tapes[pos+13993], tapes[pos+16288], tapes[pos+18583], tapes[pos+20878], tapes[pos+23173], tapes[pos+25468], tapes[pos+27763], tapes[pos+30058], tapes[pos+32353], tapes[pos+34648]};
    assign tmp_shares[3599:3584]={tapes[pos+224], tapes[pos+2519], tapes[pos+4814], tapes[pos+7109], tapes[pos+9404], tapes[pos+11699], tapes[pos+13994], tapes[pos+16289], tapes[pos+18584], tapes[pos+20879], tapes[pos+23174], tapes[pos+25469], tapes[pos+27764], tapes[pos+30059], tapes[pos+32354], tapes[pos+34649]};
    assign tmp_shares[3615:3600]={tapes[pos+225], tapes[pos+2520], tapes[pos+4815], tapes[pos+7110], tapes[pos+9405], tapes[pos+11700], tapes[pos+13995], tapes[pos+16290], tapes[pos+18585], tapes[pos+20880], tapes[pos+23175], tapes[pos+25470], tapes[pos+27765], tapes[pos+30060], tapes[pos+32355], tapes[pos+34650]};
    assign tmp_shares[3631:3616]={tapes[pos+226], tapes[pos+2521], tapes[pos+4816], tapes[pos+7111], tapes[pos+9406], tapes[pos+11701], tapes[pos+13996], tapes[pos+16291], tapes[pos+18586], tapes[pos+20881], tapes[pos+23176], tapes[pos+25471], tapes[pos+27766], tapes[pos+30061], tapes[pos+32356], tapes[pos+34651]};
    assign tmp_shares[3647:3632]={tapes[pos+227], tapes[pos+2522], tapes[pos+4817], tapes[pos+7112], tapes[pos+9407], tapes[pos+11702], tapes[pos+13997], tapes[pos+16292], tapes[pos+18587], tapes[pos+20882], tapes[pos+23177], tapes[pos+25472], tapes[pos+27767], tapes[pos+30062], tapes[pos+32357], tapes[pos+34652]};
    assign tmp_shares[3663:3648]={tapes[pos+228], tapes[pos+2523], tapes[pos+4818], tapes[pos+7113], tapes[pos+9408], tapes[pos+11703], tapes[pos+13998], tapes[pos+16293], tapes[pos+18588], tapes[pos+20883], tapes[pos+23178], tapes[pos+25473], tapes[pos+27768], tapes[pos+30063], tapes[pos+32358], tapes[pos+34653]};
    assign tmp_shares[3679:3664]={tapes[pos+229], tapes[pos+2524], tapes[pos+4819], tapes[pos+7114], tapes[pos+9409], tapes[pos+11704], tapes[pos+13999], tapes[pos+16294], tapes[pos+18589], tapes[pos+20884], tapes[pos+23179], tapes[pos+25474], tapes[pos+27769], tapes[pos+30064], tapes[pos+32359], tapes[pos+34654]};
    assign tmp_shares[3695:3680]={tapes[pos+230], tapes[pos+2525], tapes[pos+4820], tapes[pos+7115], tapes[pos+9410], tapes[pos+11705], tapes[pos+14000], tapes[pos+16295], tapes[pos+18590], tapes[pos+20885], tapes[pos+23180], tapes[pos+25475], tapes[pos+27770], tapes[pos+30065], tapes[pos+32360], tapes[pos+34655]};
    assign tmp_shares[3711:3696]={tapes[pos+231], tapes[pos+2526], tapes[pos+4821], tapes[pos+7116], tapes[pos+9411], tapes[pos+11706], tapes[pos+14001], tapes[pos+16296], tapes[pos+18591], tapes[pos+20886], tapes[pos+23181], tapes[pos+25476], tapes[pos+27771], tapes[pos+30066], tapes[pos+32361], tapes[pos+34656]};
    assign tmp_shares[3727:3712]={tapes[pos+232], tapes[pos+2527], tapes[pos+4822], tapes[pos+7117], tapes[pos+9412], tapes[pos+11707], tapes[pos+14002], tapes[pos+16297], tapes[pos+18592], tapes[pos+20887], tapes[pos+23182], tapes[pos+25477], tapes[pos+27772], tapes[pos+30067], tapes[pos+32362], tapes[pos+34657]};
    assign tmp_shares[3743:3728]={tapes[pos+233], tapes[pos+2528], tapes[pos+4823], tapes[pos+7118], tapes[pos+9413], tapes[pos+11708], tapes[pos+14003], tapes[pos+16298], tapes[pos+18593], tapes[pos+20888], tapes[pos+23183], tapes[pos+25478], tapes[pos+27773], tapes[pos+30068], tapes[pos+32363], tapes[pos+34658]};
    assign tmp_shares[3759:3744]={tapes[pos+234], tapes[pos+2529], tapes[pos+4824], tapes[pos+7119], tapes[pos+9414], tapes[pos+11709], tapes[pos+14004], tapes[pos+16299], tapes[pos+18594], tapes[pos+20889], tapes[pos+23184], tapes[pos+25479], tapes[pos+27774], tapes[pos+30069], tapes[pos+32364], tapes[pos+34659]};
    assign tmp_shares[3775:3760]={tapes[pos+235], tapes[pos+2530], tapes[pos+4825], tapes[pos+7120], tapes[pos+9415], tapes[pos+11710], tapes[pos+14005], tapes[pos+16300], tapes[pos+18595], tapes[pos+20890], tapes[pos+23185], tapes[pos+25480], tapes[pos+27775], tapes[pos+30070], tapes[pos+32365], tapes[pos+34660]};
    assign tmp_shares[3791:3776]={tapes[pos+236], tapes[pos+2531], tapes[pos+4826], tapes[pos+7121], tapes[pos+9416], tapes[pos+11711], tapes[pos+14006], tapes[pos+16301], tapes[pos+18596], tapes[pos+20891], tapes[pos+23186], tapes[pos+25481], tapes[pos+27776], tapes[pos+30071], tapes[pos+32366], tapes[pos+34661]};
    assign tmp_shares[3807:3792]={tapes[pos+237], tapes[pos+2532], tapes[pos+4827], tapes[pos+7122], tapes[pos+9417], tapes[pos+11712], tapes[pos+14007], tapes[pos+16302], tapes[pos+18597], tapes[pos+20892], tapes[pos+23187], tapes[pos+25482], tapes[pos+27777], tapes[pos+30072], tapes[pos+32367], tapes[pos+34662]};
    assign tmp_shares[3823:3808]={tapes[pos+238], tapes[pos+2533], tapes[pos+4828], tapes[pos+7123], tapes[pos+9418], tapes[pos+11713], tapes[pos+14008], tapes[pos+16303], tapes[pos+18598], tapes[pos+20893], tapes[pos+23188], tapes[pos+25483], tapes[pos+27778], tapes[pos+30073], tapes[pos+32368], tapes[pos+34663]};
    assign tmp_shares[3839:3824]={tapes[pos+239], tapes[pos+2534], tapes[pos+4829], tapes[pos+7124], tapes[pos+9419], tapes[pos+11714], tapes[pos+14009], tapes[pos+16304], tapes[pos+18599], tapes[pos+20894], tapes[pos+23189], tapes[pos+25484], tapes[pos+27779], tapes[pos+30074], tapes[pos+32369], tapes[pos+34664]};
    assign tmp_shares[3855:3840]={tapes[pos+240], tapes[pos+2535], tapes[pos+4830], tapes[pos+7125], tapes[pos+9420], tapes[pos+11715], tapes[pos+14010], tapes[pos+16305], tapes[pos+18600], tapes[pos+20895], tapes[pos+23190], tapes[pos+25485], tapes[pos+27780], tapes[pos+30075], tapes[pos+32370], tapes[pos+34665]};
    assign tmp_shares[3871:3856]={tapes[pos+241], tapes[pos+2536], tapes[pos+4831], tapes[pos+7126], tapes[pos+9421], tapes[pos+11716], tapes[pos+14011], tapes[pos+16306], tapes[pos+18601], tapes[pos+20896], tapes[pos+23191], tapes[pos+25486], tapes[pos+27781], tapes[pos+30076], tapes[pos+32371], tapes[pos+34666]};
    assign tmp_shares[3887:3872]={tapes[pos+242], tapes[pos+2537], tapes[pos+4832], tapes[pos+7127], tapes[pos+9422], tapes[pos+11717], tapes[pos+14012], tapes[pos+16307], tapes[pos+18602], tapes[pos+20897], tapes[pos+23192], tapes[pos+25487], tapes[pos+27782], tapes[pos+30077], tapes[pos+32372], tapes[pos+34667]};
    assign tmp_shares[3903:3888]={tapes[pos+243], tapes[pos+2538], tapes[pos+4833], tapes[pos+7128], tapes[pos+9423], tapes[pos+11718], tapes[pos+14013], tapes[pos+16308], tapes[pos+18603], tapes[pos+20898], tapes[pos+23193], tapes[pos+25488], tapes[pos+27783], tapes[pos+30078], tapes[pos+32373], tapes[pos+34668]};
    assign tmp_shares[3919:3904]={tapes[pos+244], tapes[pos+2539], tapes[pos+4834], tapes[pos+7129], tapes[pos+9424], tapes[pos+11719], tapes[pos+14014], tapes[pos+16309], tapes[pos+18604], tapes[pos+20899], tapes[pos+23194], tapes[pos+25489], tapes[pos+27784], tapes[pos+30079], tapes[pos+32374], tapes[pos+34669]};
    assign tmp_shares[3935:3920]={tapes[pos+245], tapes[pos+2540], tapes[pos+4835], tapes[pos+7130], tapes[pos+9425], tapes[pos+11720], tapes[pos+14015], tapes[pos+16310], tapes[pos+18605], tapes[pos+20900], tapes[pos+23195], tapes[pos+25490], tapes[pos+27785], tapes[pos+30080], tapes[pos+32375], tapes[pos+34670]};
    assign tmp_shares[3951:3936]={tapes[pos+246], tapes[pos+2541], tapes[pos+4836], tapes[pos+7131], tapes[pos+9426], tapes[pos+11721], tapes[pos+14016], tapes[pos+16311], tapes[pos+18606], tapes[pos+20901], tapes[pos+23196], tapes[pos+25491], tapes[pos+27786], tapes[pos+30081], tapes[pos+32376], tapes[pos+34671]};
    assign tmp_shares[3967:3952]={tapes[pos+247], tapes[pos+2542], tapes[pos+4837], tapes[pos+7132], tapes[pos+9427], tapes[pos+11722], tapes[pos+14017], tapes[pos+16312], tapes[pos+18607], tapes[pos+20902], tapes[pos+23197], tapes[pos+25492], tapes[pos+27787], tapes[pos+30082], tapes[pos+32377], tapes[pos+34672]};
    assign tmp_shares[3983:3968]={tapes[pos+248], tapes[pos+2543], tapes[pos+4838], tapes[pos+7133], tapes[pos+9428], tapes[pos+11723], tapes[pos+14018], tapes[pos+16313], tapes[pos+18608], tapes[pos+20903], tapes[pos+23198], tapes[pos+25493], tapes[pos+27788], tapes[pos+30083], tapes[pos+32378], tapes[pos+34673]};
    assign tmp_shares[3999:3984]={tapes[pos+249], tapes[pos+2544], tapes[pos+4839], tapes[pos+7134], tapes[pos+9429], tapes[pos+11724], tapes[pos+14019], tapes[pos+16314], tapes[pos+18609], tapes[pos+20904], tapes[pos+23199], tapes[pos+25494], tapes[pos+27789], tapes[pos+30084], tapes[pos+32379], tapes[pos+34674]};
    assign tmp_shares[4015:4000]={tapes[pos+250], tapes[pos+2545], tapes[pos+4840], tapes[pos+7135], tapes[pos+9430], tapes[pos+11725], tapes[pos+14020], tapes[pos+16315], tapes[pos+18610], tapes[pos+20905], tapes[pos+23200], tapes[pos+25495], tapes[pos+27790], tapes[pos+30085], tapes[pos+32380], tapes[pos+34675]};
    assign tmp_shares[4031:4016]={tapes[pos+251], tapes[pos+2546], tapes[pos+4841], tapes[pos+7136], tapes[pos+9431], tapes[pos+11726], tapes[pos+14021], tapes[pos+16316], tapes[pos+18611], tapes[pos+20906], tapes[pos+23201], tapes[pos+25496], tapes[pos+27791], tapes[pos+30086], tapes[pos+32381], tapes[pos+34676]};
    assign tmp_shares[4047:4032]={tapes[pos+252], tapes[pos+2547], tapes[pos+4842], tapes[pos+7137], tapes[pos+9432], tapes[pos+11727], tapes[pos+14022], tapes[pos+16317], tapes[pos+18612], tapes[pos+20907], tapes[pos+23202], tapes[pos+25497], tapes[pos+27792], tapes[pos+30087], tapes[pos+32382], tapes[pos+34677]};
    assign tmp_shares[4063:4048]={tapes[pos+253], tapes[pos+2548], tapes[pos+4843], tapes[pos+7138], tapes[pos+9433], tapes[pos+11728], tapes[pos+14023], tapes[pos+16318], tapes[pos+18613], tapes[pos+20908], tapes[pos+23203], tapes[pos+25498], tapes[pos+27793], tapes[pos+30088], tapes[pos+32383], tapes[pos+34678]};
    assign tmp_shares[4079:4064]={tapes[pos+254], tapes[pos+2549], tapes[pos+4844], tapes[pos+7139], tapes[pos+9434], tapes[pos+11729], tapes[pos+14024], tapes[pos+16319], tapes[pos+18614], tapes[pos+20909], tapes[pos+23204], tapes[pos+25499], tapes[pos+27794], tapes[pos+30089], tapes[pos+32384], tapes[pos+34679]};
    
    

endmodule


module mpc_AND3(//this module is for signature generation
    input a,
    input b,
    input [15:0] mask_a,
    input [15:0] mask_b,
    input [`tapesLength-1:0] tapes,
    input [`msgsLength-1:0] msgs,
    input [10:0] tapesPos,
    input [10:0] msgsPos,
    
    output [`msgsLength-1:0] updated_msgs,
    output c
    );
    
    wire [15:0] and_helper;
    wire [15:0] s_shares;
    wire [15:0] extended_a;
    wire [15:0] extended_b;
    wire [`one_msgsLength-1:0] result_helper0;
    wire parity_s_shares;
    wire [`one_msgsLength-1:0] temp0, temp1, temp2, temp3, temp4, temp5, temp6, temp7, temp8, temp9, temp10, temp11, temp12, temp13, temp14, temp15;
    
    
    assign and_helper={tapes[tapesPos],tapes[tapesPos+2295],tapes[tapesPos+4590],tapes[tapesPos+6885],tapes[tapesPos+9180],tapes[tapesPos+11475],tapes[tapesPos+13770],tapes[tapesPos+16065],tapes[tapesPos+18360],tapes[tapesPos+20655],tapes[tapesPos+22950],tapes[tapesPos+25245],tapes[tapesPos+27540],tapes[tapesPos+29835],tapes[tapesPos+32130],tapes[tapesPos+34425]};
    assign extended_a={a, a, a, a, a, a, a, a, a, a, a, a, a, a, a, a};
    assign extended_b={b, b, b, b, b, b, b, b, b, b, b, b, b, b, b};
    assign s_shares=(extended_a & mask_b) ^ (extended_b & mask_a) ^ and_helper;
    assign parity_s_shares=s_shares[0] ^  s_shares[1] ^  s_shares[2] ^  s_shares[3] ^  s_shares[4] ^  s_shares[5] ^  s_shares[6] ^  s_shares[7] ^  s_shares[8] ^  s_shares[9] ^  s_shares[10] ^  s_shares[11] ^  s_shares[12] ^  s_shares[13] ^  s_shares[14] ^  s_shares[15];
    assign c=parity_s_shares ^ (a & b);
    
    assign result_helper0=1275'b1<<(msgsPos);

    
    assign temp0=(s_shares[0]==1)? (msgs[1274:0] | result_helper0) : (msgs[1274:0] & ~result_helper0);
    assign temp1=(s_shares[1]==1)? (msgs[2549:1275] | result_helper0) : (msgs[2549:1275] & ~result_helper0);
    assign temp2=(s_shares[2]==1)? (msgs[3824:2550] | result_helper0) : (msgs[3824:2550] & ~result_helper0);
    assign temp3=(s_shares[3]==1)? (msgs[5099:3825] | result_helper0) : (msgs[5099:3825] & ~result_helper0);
    assign temp4=(s_shares[4]==1)? (msgs[6374:5100] | result_helper0) : (msgs[6374:5100] & ~result_helper0);
    assign temp5=(s_shares[5]==1)? (msgs[7649:6375] | result_helper0) : (msgs[7649:6375] & ~result_helper0);
    assign temp6=(s_shares[6]==1)? (msgs[8924:7650] | result_helper0) : (msgs[8924:7650] & ~result_helper0);
    assign temp7=(s_shares[7]==1)? (msgs[10199:8925] | result_helper0) : (msgs[10199:8925] & ~result_helper0);
    assign temp8=(s_shares[8]==1)? (msgs[11474:10200] | result_helper0) : (msgs[11474:10200] & ~result_helper0);
    assign temp9=(s_shares[9]==1)? (msgs[12749:11475] | result_helper0) : (msgs[12749:11475] & ~result_helper0);
    assign temp10=(s_shares[10]==1)? (msgs[14024:12750] | result_helper0) : (msgs[14024:12750] & ~result_helper0);
    assign temp11=(s_shares[11]==1)? (msgs[16574:15300] | result_helper0) : (msgs[16574:15300] & ~result_helper0);
    assign temp12=(s_shares[12]==1)? (msgs[17849:16575] | result_helper0) : (msgs[17849:16575] & ~result_helper0);
    assign temp13=(s_shares[13]==1)? (msgs[17849:16575] | result_helper0) : (msgs[17849:16575] & ~result_helper0);
    assign temp14=(s_shares[14]==1)? (msgs[19124:17850] | result_helper0) : (msgs[19124:17850] & ~result_helper0);
    assign temp15=(s_shares[15]==1)? (msgs[20399:19125] | result_helper0) : (msgs[20399:19125] & ~result_helper0);
    
    assign updated_msgs[1274:0]=temp0;//
    assign updated_msgs[2549:1275]=temp1;//
    assign updated_msgs[3824:2550]=temp2;//
    assign updated_msgs[5099:3825]=temp3;//
    assign updated_msgs[6374:5100]=temp4;//
    assign updated_msgs[7649:6375]=temp5;//
    assign updated_msgs[8924:7650]=temp6;//
    assign updated_msgs[10199:8925]=temp7;
    assign updated_msgs[11474:10200]=temp8;
    assign updated_msgs[12749:11475]=temp9;
    assign updated_msgs[14024:12750]=temp10;
    assign updated_msgs[15299:14025]=temp11;
    assign updated_msgs[16574:15300]=temp12;
    assign updated_msgs[17849:16575]=temp13;
    assign updated_msgs[19124:17850]=temp14;
    assign updated_msgs[20399:19125]=temp15;//
    
endmodule


module mpc_AND33(
    input a,
    input b,
    input c,
    input [15:0] mask_a,
    input [15:0] mask_b,
    input [15:0] mask_c,
    input [`tapesLength-1:0] tapes,
    input [`msgsLength-1:0] msgs,
    input [10:0] tapesPos,
    input [10:0] msgsPos,
    
    output [`msgsLength-1:0] updated_msgs,
    output ab,
    output bc,
    output ca
);
    wire [`msgsLength-1:0] FirstTime_msgs_Result, SecondTime_msgs_Result, ThirdTime_msgs_Result;

    wire ab_temp, bc_temp, ca_temp;
    
    
    mpc_AND3 FirstTime(a, b, mask_a, mask_b, tapes, msgs, tapesPos, msgsPos, FirstTime_msgs_Result, ab_temp);
    
    
    mpc_AND3 SecondTime(b, c, mask_b, mask_c, tapes, FirstTime_msgs_Result, tapesPos+1, msgsPos+1, SecondTime_msgs_Result, bc_temp);
    
    
    mpc_AND3 ThirdTime(c, a, mask_c, mask_a, tapes, SecondTime_msgs_Result, tapesPos+2, msgsPos+2, ThirdTime_msgs_Result, ca_temp);
    
    
    assign ab=ab_temp;
    assign bc=bc_temp;
    assign ca=ca_temp;
    assign updated_msgs=ThirdTime_msgs_Result;
endmodule






module mpc_sbox3(
    input clk,
    input rst,
    input start,
    input [254:0] state,
    input [`state_mask_length-1:0] state_mask,
    input [`tapesLength-1:0] tapes,
    input [`msgsLength-1:0] msgs,
    input [10:0] tapesPos,
    input [10:0] msgsPos,
    
    output [254:0] updated_state,
    output [`msgsLength-1:0] updated_msgs,
    output stop
);
    
    wire a, b, c, ab, bc, ca;
    wire [15:0] mask_a, mask_b, mask_c;
    wire [`msgsLength-1:0] new_msgs; 
    wire state_updated1, state_updated2, state_updated3;
    reg [7:0] i;
    reg [`msgsLength-1:0] msgs_reg;
    reg [254:0] state_reg;
    reg [10:0] tapesPos_reg, msgsPos_reg;
    reg stop_reg;
    reg [1:0] ControlState;
    
    
    assign a=state_reg[i+2];
    assign mask_a={state_mask[(i+2)*16+15], state_mask[(i+2)*16+14], state_mask[(i+2)*16+13], state_mask[(i+2)*16+12], state_mask[(i+2)*16+11], state_mask[(i+2)*16+10], state_mask[(i+2)*16+9], state_mask[(i+2)*16+8], state_mask[(i+2)*16+7], state_mask[(i+2)*16+6], state_mask[(i+2)*16+5], state_mask[(i+2)*16+4], state_mask[(i+2)*16+3], state_mask[(i+2)*16+2], state_mask[(i+2)*16+1], state_mask[(i+2)*16] };
    
    assign b=state_reg[i+1];
    assign mask_b={state_mask[(i+1)*16+15], state_mask[(i+1)*16+14], state_mask[(i+1)*16+13], state_mask[(i+1)*16+12], state_mask[(i+1)*16+11], state_mask[(i+1)*16+10], state_mask[(i+1)*16+9], state_mask[(i+1)*16+8], state_mask[(i+1)*16+7], state_mask[(i+1)*16+6], state_mask[(i+1)*16+5], state_mask[(i+1)*16+4], state_mask[(i+1)*16+3], state_mask[(i+1)*16+2], state_mask[(i+1)*16+1], state_mask[(i+1)*16] };
    
    assign c=state_reg[i];
    assign mask_c={state_mask[(i)*16], state_mask[(i)*16+1], state_mask[(i)*16+2], state_mask[(i)*16+3], state_mask[(i)*16+4], state_mask[(i)*16+5], state_mask[(i)*16+6], state_mask[(i)*16+7], state_mask[(i)*16+8], state_mask[(i)*16+9], state_mask[(i)*16+10], state_mask[(i)*16+11], state_mask[(i)*16+12], state_mask[(i)*16+13], state_mask[(i)*16+14], state_mask[(i)*16+15]};
    
    mpc_AND33 Three3TimesAND(a, b, c, mask_a, mask_b, mask_c, tapes, msgs_reg, tapesPos_reg, msgsPos_reg, new_msgs, ab, bc, ca);
    
    assign state_updated1=a ^ bc;
    assign state_updated2=a ^ b ^ ca;
    assign state_updated3=a ^ b ^ c ^ ab;

    //control
    always@(posedge clk or negedge rst)
    begin
        if(!rst)
            begin
                ControlState<=2'b00;
            end
        else
            begin
                if(ControlState==2'b00)
                    begin
                        stop_reg<=0;
                        if(start)
                            begin
                                tapesPos_reg<=tapesPos;
                                msgsPos_reg<=msgsPos;
                                msgs_reg<=msgs;
                                state_reg<=state;
                                i<=0;
                                ControlState<=2'b01;
                            end
                    end
                    
                else if(ControlState==2'b01)
                    begin
                        if(i!=252)
                            begin
                                i<=i+3;
                                msgs_reg<=new_msgs;
                                tapesPos_reg<=tapesPos_reg+3;
                                msgsPos_reg<=msgsPos_reg+3;
                                
                                state_reg[i+2]<=state_updated1;
                                state_reg[i+1]<=state_updated2;
                                state_reg[i]<=state_updated3;
                            end
                        else
                            begin
                                ControlState<=2'b10;
                            end
                    end
                
                else if(ControlState==2'b10)
                    begin
                        i<=252;
                        ControlState<=2'b11;
                        state_reg[i+2]<=state_updated1;
                        state_reg[i+1]<=state_updated2;
                        state_reg[i]<=state_updated3;
                        stop_reg<=1;
                    end
                else if(ControlState==2'b11)
                    begin
                        stop_reg<=1;
                        ControlState<=2'b00;
                    end
            end
    end

    //output
    assign stop=stop_reg;
    assign updated_state=state_reg;
    assign updated_msgs=msgs_reg;
endmodule





module mpc_simulate(
    input clk,
    input rst,
    input start,
    input [254:0] masked_key,
    input [254: 0] C,
    input [254:0] p,
    input [`tapesLength-1:0] tapes,
    input [`msgsLength-1:0] msgs,
    
    output[`msgsLength-1:0] updated_msgs,
    output stop
);
    
    wire [254:0] initial_whitening_round_key;
    wire [254:0] initial_whitening_state;
    wire [254:0] updated_state;
    wire [`msgsLength-1:0] new_msgs;
    wire inside_stop;
    wire [254:0] Matrix_mul_Result;
    wire [254:0] Add_Round_Constant_Result;
    wire [254:0] round_key;
    wire [254:0] Add_Round_Key_Result;
    wire [`state_mask_length-1:0] tmp_shares_wire;
    
    reg [1:0] round;
    reg [254:0] state;
    //reg [`state_mask_length-1:0] tmp_shares;
    //reg [`tapesLength-1:0] tapes_reg;
    reg [`msgsLength-1:0] msgs_reg;
    reg [10:0] tapesPos_reg;
    reg [10:0] msgsPos_reg;
    reg stop_reg, start_reg;
    reg [3:0] ControlState;
    
    //---------------------------Initial Whitening------------------------------
    compute_whitening_key CWK(masked_key, initial_whitening_round_key);
    assign initial_whitening_state=p^initial_whitening_round_key;
    
    
    //---------------------------LowMC Rounds with mpc_sbox3 as sbox layer-------------------------------
    tapes2tmp_shares T2T(tapes, tapesPos_reg, tmp_shares_wire);
    mpc_sbox3 SBOX(clk, rst, start_reg, state, tmp_shares_wire, tapes, msgs_reg, tapesPos_reg, msgsPos_reg, updated_state, new_msgs, inside_stop);
    Matrix_Multiplication MUL(updated_state, round, Matrix_mul_Result);
    Add_Constant ADDC(Matrix_mul_Result, round, Add_Round_Constant_Result);
    Key_Expansion EXP(masked_key, round, round_key);
    assign Add_Round_Key_Result=round_key ^ Add_Round_Constant_Result;
    
    
    //control
    always@(posedge clk or negedge rst)
    begin
        if(!rst)
            begin
                ControlState<=0;
                start_reg<=0;
            end
        else
            begin
            
            
                if(ControlState==0)
                    begin
                        stop_reg<=0;
                        if(start)
                            begin
                                msgs_reg<=msgs;
                                state<=initial_whitening_state;
                                round<=2'b00;
                                tapesPos_reg<=11'b0;
                                msgsPos_reg<=11'b0;
                                start_reg<=0;
                                ControlState<=1;
                            end
                    end
                    
                else if(ControlState==1)
                    begin
                        start_reg<=1;
                        if(inside_stop)
                            begin
                                start_reg<=0;
                                ControlState<=2;
                            end
                    end
                    
                else if(ControlState==2)
                    begin
                        msgs_reg<=new_msgs;
                        state<=updated_state;
                        round<=2'b01;
                        tapesPos_reg<=2*255;
                        msgsPos_reg<=255;
                        ControlState<=3;
                    end
                    
                else if(ControlState==3)
                    begin
                        start_reg<=1;
                        if(inside_stop)
                            begin
                                start_reg<=0;
                                ControlState<=4;
                            end
                    end
                    
                else if(ControlState==4)
                    begin
                        msgs_reg<=new_msgs;
                        state<=updated_state;
                        round<=2'b10;
                        tapesPos_reg<=4*255;
                        msgsPos_reg<=2*255;
                        ControlState<=5;
                    end
                    
                else if(ControlState==5)
                    begin
                        start_reg<=1;
                        if(inside_stop)
                            begin
                                start_reg<=0;
                                ControlState<=6;
                            end
                    end
                    
                else if(ControlState==6)
                    begin
                        msgs_reg<=new_msgs;
                        state<=updated_state;
                        round<=2'b11;
                        tapesPos_reg<=6*255;
                        msgsPos_reg<=3*255;
                        ControlState<=7;
                    end
                    
                else if(ControlState==7)
                    begin
                        start_reg<=1;
                        if(inside_stop)
                            begin
                                stop_reg<=1;
                                start_reg<=0;
                                ControlState<=0;
                            end
                    end
                    
                    
            end
    end
    
    
    assign stop=stop_reg;
    assign updated_msgs=new_msgs;
    //assign inside=inside_stop;
    //assign state_out=ControlState;
    //assign inside_start=start_reg;
endmodule
    
    
    
    