`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/02 23:39:15
// Design Name: 
// Module Name: simulate_part1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module simulate_part1(
    input [254:0] Lambda_mpc,
    input [7:0] a,
    
    output [7:0] part1
    );
    
    assign part1[0]=((a[5]) & Lambda_mpc[1] ^ Lambda_mpc[5]) ^ ((a[6]) & Lambda_mpc[3] ^ Lambda_mpc[5]) ^ (a[5] & a[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[6]) ^ (a[5] & a[6] & a[7]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[159] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[143] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
    assign part1[1]=(a[7]) ^ ((a[6]) & Lambda_mpc[0] ^ Lambda_mpc[2]) ^ ((a[7]) & Lambda_mpc[1] ^ Lambda_mpc[2]) ^ (a[6] & a[7]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[6]) ^ (a[5] & a[6] & a[7]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[14]) ^ (a[4] & a[5] & a[6] & a[7]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[191] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[135] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
    assign part1[2]=(a[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[6]) ^ (a[5] & a[6] & a[7]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[14]) ^ (a[4] & a[5] & a[6] & a[7]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[62]) ^ (a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[126]) ^ (a[1] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[159] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[143] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[135] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
    assign part1[3]=(a[6]) ^ ((a[6]) & Lambda_mpc[0] ^ Lambda_mpc[2]) ^ ((a[7]) & Lambda_mpc[1] ^ Lambda_mpc[2]) ^ (a[6] & a[7]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[6]) ^ (a[5] & a[6] & a[7]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[14]) ^ (a[4] & a[5] & a[6] & a[7]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[131] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
    assign part1[4]=(a[6]) ^ ((a[5]) & Lambda_mpc[1] ^ Lambda_mpc[5]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[14]) ^ (a[4] & a[5] & a[6] & a[7]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[62]) ^ (a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[191] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[159] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[143] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[135] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[131] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]);
    assign part1[5]=(a[7]) ^ ((a[6]) & Lambda_mpc[0] ^ Lambda_mpc[2]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[6]) ^ (a[5] & a[6] & a[7]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[126]) ^ (a[1] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[191] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[143] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[129] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
    assign part1[6]=(a[7]) ^ ((a[6]) & Lambda_mpc[0] ^ Lambda_mpc[2]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[6]) & Lambda_mpc[4] ^ Lambda_mpc[6]) ^ ((a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[6]) ^ (a[5] & a[6] & a[7]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[5]) & Lambda_mpc[10] ^ Lambda_mpc[14]) ^ ((a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[14]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[14]) ^ (a[4] & a[5] & a[6] & a[7]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[30]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[30]) ^ (a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[62]) ^ (a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[126]) ^ (a[1] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[195] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[199] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[191] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[147] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[151] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[143] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
    assign part1[7]=(a[6]) ^ ((a[6]) & Lambda_mpc[0] ^ Lambda_mpc[2]) ^ ((a[7]) & Lambda_mpc[1] ^ Lambda_mpc[2]) ^ (a[6] & a[7]) ^ ((a[5]) & Lambda_mpc[2] ^ Lambda_mpc[6]) ^ ((a[7]) & Lambda_mpc[5] ^ Lambda_mpc[6]) ^ ((a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[6]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[4]) & Lambda_mpc[6] ^ Lambda_mpc[14]) ^ ((a[6]) & Lambda_mpc[12] ^ Lambda_mpc[14]) ^ ((a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[14]) ^ ((a[7]) & Lambda_mpc[13] ^ Lambda_mpc[14]) ^ ((a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[14]) ^ ((a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[14]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[14]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[30]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[30]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[7]) & Lambda_mpc[29] ^ Lambda_mpc[30]) ^ ((a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[30]) ^ ((a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[30]) ^ ((a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[30]) ^ ((a[3]) & Lambda_mpc[14] ^ Lambda_mpc[30]) ^ ((a[4]) & Lambda_mpc[22] ^ Lambda_mpc[30]) ^ ((a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[30]) ^ ((a[5]) & Lambda_mpc[26] ^ Lambda_mpc[30]) ^ ((a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[30]) ^ ((a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[30]) ^ ((a[6]) & Lambda_mpc[28] ^ Lambda_mpc[30]) ^ ((a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[30]) ^ ((a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[30]) ^ ((a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[30]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[30]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[30]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[30]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[2]) & Lambda_mpc[30] ^ Lambda_mpc[62]) ^ ((a[3]) & Lambda_mpc[46] ^ Lambda_mpc[62]) ^ ((a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[62]) ^ ((a[4]) & Lambda_mpc[54] ^ Lambda_mpc[62]) ^ ((a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[62]) ^ ((a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[62]) ^ ((a[5]) & Lambda_mpc[58] ^ Lambda_mpc[62]) ^ ((a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[62]) ^ ((a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[62]) ^ ((a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[62]) ^ ((a[6]) & Lambda_mpc[60] ^ Lambda_mpc[62]) ^ ((a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[62]) ^ ((a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[62]) ^ ((a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[62]) ^ ((a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[62]) ^ ((a[7]) & Lambda_mpc[61] ^ Lambda_mpc[62]) ^ ((a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[62]) ^ ((a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[62]) ^ ((a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[62]) ^ ((a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[62]) ^ ((a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[62]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[62]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[62]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[62]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[62]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[62]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[62]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[62]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[62]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[62]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[62]) ^ (a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[1]) & Lambda_mpc[62] ^ Lambda_mpc[126]) ^ ((a[2]) & Lambda_mpc[94] ^ Lambda_mpc[126]) ^ ((a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[126]) ^ ((a[3]) & Lambda_mpc[110] ^ Lambda_mpc[126]) ^ ((a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[126]) ^ ((a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[126]) ^ ((a[4]) & Lambda_mpc[118] ^ Lambda_mpc[126]) ^ ((a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[126]) ^ ((a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[126]) ^ ((a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[126]) ^ ((a[5]) & Lambda_mpc[122] ^ Lambda_mpc[126]) ^ ((a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[126]) ^ ((a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[126]) ^ ((a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[126]) ^ ((a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[126]) ^ ((a[6]) & Lambda_mpc[124] ^ Lambda_mpc[126]) ^ ((a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[126]) ^ ((a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[126]) ^ ((a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[126]) ^ ((a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[126]) ^ ((a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[126]) ^ ((a[7]) & Lambda_mpc[125] ^ Lambda_mpc[126]) ^ ((a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[126]) ^ ((a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[126]) ^ ((a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[126]) ^ ((a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[126]) ^ ((a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[126]) ^ ((a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[126]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[126]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[126]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[126]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[19] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[67] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[3] ^ Lambda_mpc[126]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[126]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[126]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[23] ^ Lambda_mpc[126]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[71] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[7] ^ Lambda_mpc[126]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[126]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[126]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[126]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[15] ^ Lambda_mpc[126]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[126]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[126]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[63] ^ Lambda_mpc[126]) ^ (a[1] & a[2] & a[3] & a[4] & a[5] & a[6] & a[7]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[211] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6] & a[7]) & Lambda_mpc[83] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[215] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6] & a[7]) & Lambda_mpc[87] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[207] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[79] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[4] & a[6] & a[7]) & Lambda_mpc[243] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6] & a[7]) & Lambda_mpc[115] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[179] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6] & a[7]) & Lambda_mpc[51] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[227] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[99] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[163] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6] & a[7]) & Lambda_mpc[35] ^ Lambda_mpc[254]) ^ ((a[5] & a[6] & a[7]) & Lambda_mpc[247] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6] & a[7]) & Lambda_mpc[119] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[183] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6] & a[7]) & Lambda_mpc[55] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[231] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[103] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[167] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6] & a[7]) & Lambda_mpc[39] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[239] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[111] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[175] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[47] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[223] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[95] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[159] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6] & a[7]) & Lambda_mpc[31] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[6] & a[7]) & Lambda_mpc[251] ^ Lambda_mpc[254]) ^ ((a[0] & a[6] & a[7]) & Lambda_mpc[123] ^ Lambda_mpc[254]) ^ ((a[1] & a[6] & a[7]) & Lambda_mpc[187] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6] & a[7]) & Lambda_mpc[59] ^ Lambda_mpc[254]) ^ ((a[2] & a[6] & a[7]) & Lambda_mpc[219] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6] & a[7]) & Lambda_mpc[91] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[155] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6] & a[7]) & Lambda_mpc[27] ^ Lambda_mpc[254]) ^ ((a[3] & a[6] & a[7]) & Lambda_mpc[235] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6] & a[7]) & Lambda_mpc[107] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[171] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6] & a[7]) & Lambda_mpc[43] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[203] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[75] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[139] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6] & a[7]) & Lambda_mpc[11] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[7]) & Lambda_mpc[253] ^ Lambda_mpc[254]) ^ ((a[0] & a[7]) & Lambda_mpc[125] ^ Lambda_mpc[254]) ^ ((a[1] & a[7]) & Lambda_mpc[189] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[7]) & Lambda_mpc[61] ^ Lambda_mpc[254]) ^ ((a[2] & a[7]) & Lambda_mpc[221] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[7]) & Lambda_mpc[93] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[7]) & Lambda_mpc[157] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[7]) & Lambda_mpc[29] ^ Lambda_mpc[254]) ^ ((a[3] & a[7]) & Lambda_mpc[237] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[7]) & Lambda_mpc[109] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[7]) & Lambda_mpc[173] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[7]) & Lambda_mpc[45] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[7]) & Lambda_mpc[205] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[7]) & Lambda_mpc[77] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[141] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[7]) & Lambda_mpc[13] ^ Lambda_mpc[254]) ^ ((a[4] & a[7]) & Lambda_mpc[245] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[7]) & Lambda_mpc[117] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[7]) & Lambda_mpc[181] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[7]) & Lambda_mpc[53] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[7]) & Lambda_mpc[213] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[7]) & Lambda_mpc[85] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[149] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[7]) & Lambda_mpc[21] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[7]) & Lambda_mpc[229] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[7]) & Lambda_mpc[101] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[165] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[7]) & Lambda_mpc[37] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[197] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[69] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[133] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[7]) & Lambda_mpc[5] ^ Lambda_mpc[254]) ^ ((a[5] & a[7]) & Lambda_mpc[249] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[7]) & Lambda_mpc[121] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[7]) & Lambda_mpc[185] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[7]) & Lambda_mpc[57] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[7]) & Lambda_mpc[217] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[7]) & Lambda_mpc[89] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[153] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[7]) & Lambda_mpc[25] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[7]) & Lambda_mpc[233] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[7]) & Lambda_mpc[105] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[169] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[7]) & Lambda_mpc[41] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[201] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[73] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[137] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[7]) & Lambda_mpc[9] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[7]) & Lambda_mpc[241] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[7]) & Lambda_mpc[113] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[177] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[7]) & Lambda_mpc[49] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[209] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[81] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[145] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[7]) & Lambda_mpc[17] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[225] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[97] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[161] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[33] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[193] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[65] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[129] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[7]) & Lambda_mpc[1] ^ Lambda_mpc[254]) ^ ((a[0]) & Lambda_mpc[126] ^ Lambda_mpc[254]) ^ ((a[1]) & Lambda_mpc[190] ^ Lambda_mpc[254]) ^ ((a[0] & a[1]) & Lambda_mpc[62] ^ Lambda_mpc[254]) ^ ((a[2]) & Lambda_mpc[222] ^ Lambda_mpc[254]) ^ ((a[0] & a[2]) & Lambda_mpc[94] ^ Lambda_mpc[254]) ^ ((a[1] & a[2]) & Lambda_mpc[158] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2]) & Lambda_mpc[30] ^ Lambda_mpc[254]) ^ ((a[3]) & Lambda_mpc[238] ^ Lambda_mpc[254]) ^ ((a[0] & a[3]) & Lambda_mpc[110] ^ Lambda_mpc[254]) ^ ((a[1] & a[3]) & Lambda_mpc[174] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3]) & Lambda_mpc[46] ^ Lambda_mpc[254]) ^ ((a[2] & a[3]) & Lambda_mpc[206] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3]) & Lambda_mpc[78] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3]) & Lambda_mpc[142] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3]) & Lambda_mpc[14] ^ Lambda_mpc[254]) ^ ((a[4]) & Lambda_mpc[246] ^ Lambda_mpc[254]) ^ ((a[0] & a[4]) & Lambda_mpc[118] ^ Lambda_mpc[254]) ^ ((a[1] & a[4]) & Lambda_mpc[182] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4]) & Lambda_mpc[54] ^ Lambda_mpc[254]) ^ ((a[2] & a[4]) & Lambda_mpc[214] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4]) & Lambda_mpc[86] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4]) & Lambda_mpc[150] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4]) & Lambda_mpc[22] ^ Lambda_mpc[254]) ^ ((a[3] & a[4]) & Lambda_mpc[230] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4]) & Lambda_mpc[102] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4]) & Lambda_mpc[166] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4]) & Lambda_mpc[38] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4]) & Lambda_mpc[198] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4]) & Lambda_mpc[70] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[134] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4]) & Lambda_mpc[6] ^ Lambda_mpc[254]) ^ ((a[5]) & Lambda_mpc[250] ^ Lambda_mpc[254]) ^ ((a[0] & a[5]) & Lambda_mpc[122] ^ Lambda_mpc[254]) ^ ((a[1] & a[5]) & Lambda_mpc[186] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5]) & Lambda_mpc[58] ^ Lambda_mpc[254]) ^ ((a[2] & a[5]) & Lambda_mpc[218] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5]) & Lambda_mpc[90] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5]) & Lambda_mpc[154] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5]) & Lambda_mpc[26] ^ Lambda_mpc[254]) ^ ((a[3] & a[5]) & Lambda_mpc[234] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5]) & Lambda_mpc[106] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5]) & Lambda_mpc[170] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5]) & Lambda_mpc[42] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5]) & Lambda_mpc[202] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5]) & Lambda_mpc[74] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[138] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5]) & Lambda_mpc[10] ^ Lambda_mpc[254]) ^ ((a[4] & a[5]) & Lambda_mpc[242] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5]) & Lambda_mpc[114] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5]) & Lambda_mpc[178] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5]) & Lambda_mpc[50] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5]) & Lambda_mpc[210] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5]) & Lambda_mpc[82] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[146] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5]) & Lambda_mpc[18] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5]) & Lambda_mpc[226] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5]) & Lambda_mpc[98] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[162] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5]) & Lambda_mpc[34] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[194] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[66] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[130] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5]) & Lambda_mpc[2] ^ Lambda_mpc[254]) ^ ((a[6]) & Lambda_mpc[252] ^ Lambda_mpc[254]) ^ ((a[0] & a[6]) & Lambda_mpc[124] ^ Lambda_mpc[254]) ^ ((a[1] & a[6]) & Lambda_mpc[188] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[6]) & Lambda_mpc[60] ^ Lambda_mpc[254]) ^ ((a[2] & a[6]) & Lambda_mpc[220] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[6]) & Lambda_mpc[92] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[6]) & Lambda_mpc[156] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[6]) & Lambda_mpc[28] ^ Lambda_mpc[254]) ^ ((a[3] & a[6]) & Lambda_mpc[236] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[6]) & Lambda_mpc[108] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[6]) & Lambda_mpc[172] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[6]) & Lambda_mpc[44] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[6]) & Lambda_mpc[204] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[6]) & Lambda_mpc[76] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[140] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[6]) & Lambda_mpc[12] ^ Lambda_mpc[254]) ^ ((a[4] & a[6]) & Lambda_mpc[244] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[6]) & Lambda_mpc[116] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[6]) & Lambda_mpc[180] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[6]) & Lambda_mpc[52] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[6]) & Lambda_mpc[212] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[6]) & Lambda_mpc[84] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[148] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[6]) & Lambda_mpc[20] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[6]) & Lambda_mpc[228] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[6]) & Lambda_mpc[100] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[164] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[6]) & Lambda_mpc[36] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[196] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[68] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[132] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[6]) & Lambda_mpc[4] ^ Lambda_mpc[254]) ^ ((a[5] & a[6]) & Lambda_mpc[248] ^ Lambda_mpc[254]) ^ ((a[0] & a[5] & a[6]) & Lambda_mpc[120] ^ Lambda_mpc[254]) ^ ((a[1] & a[5] & a[6]) & Lambda_mpc[184] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[5] & a[6]) & Lambda_mpc[56] ^ Lambda_mpc[254]) ^ ((a[2] & a[5] & a[6]) & Lambda_mpc[216] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[5] & a[6]) & Lambda_mpc[88] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[152] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[5] & a[6]) & Lambda_mpc[24] ^ Lambda_mpc[254]) ^ ((a[3] & a[5] & a[6]) & Lambda_mpc[232] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[5] & a[6]) & Lambda_mpc[104] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[168] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[5] & a[6]) & Lambda_mpc[40] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[200] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[72] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[136] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[5] & a[6]) & Lambda_mpc[8] ^ Lambda_mpc[254]) ^ ((a[4] & a[5] & a[6]) & Lambda_mpc[240] ^ Lambda_mpc[254]) ^ ((a[0] & a[4] & a[5] & a[6]) & Lambda_mpc[112] ^ Lambda_mpc[254]) ^ ((a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[176] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[4] & a[5] & a[6]) & Lambda_mpc[48] ^ Lambda_mpc[254]) ^ ((a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[208] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[80] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[144] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[4] & a[5] & a[6]) & Lambda_mpc[16] ^ Lambda_mpc[254]) ^ ((a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[224] ^ Lambda_mpc[254]) ^ ((a[0] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[96] ^ Lambda_mpc[254]) ^ ((a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[160] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[32] ^ Lambda_mpc[254]) ^ ((a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[192] ^ Lambda_mpc[254]) ^ ((a[0] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[64] ^ Lambda_mpc[254]) ^ ((a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[128] ^ Lambda_mpc[254]) ^ ((a[0] & a[1] & a[2] & a[3] & a[4] & a[5] & a[6]) & Lambda_mpc[0] ^ Lambda_mpc[254]);
endmodule



